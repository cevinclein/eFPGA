VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO LUT4AB
  CLASS BLOCK ;
  FOREIGN LUT4AB ;
  ORIGIN 0.000 0.000 ;
  SIZE 225.000 BY 225.000 ;
  PIN Ci
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 0.800 ;
    END
  END Ci
  PIN Co
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 170.750 224.200 171.030 225.000 ;
    END
  END Co
  PIN E1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 91.160 225.000 91.760 ;
    END
  END E1BEG[0]
  PIN E1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 92.520 225.000 93.120 ;
    END
  END E1BEG[1]
  PIN E1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 93.880 225.000 94.480 ;
    END
  END E1BEG[2]
  PIN E1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 95.240 225.000 95.840 ;
    END
  END E1BEG[3]
  PIN E1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 0.800 91.760 ;
    END
  END E1END[0]
  PIN E1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 0.800 93.120 ;
    END
  END E1END[1]
  PIN E1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 0.800 94.480 ;
    END
  END E1END[2]
  PIN E1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 0.800 95.840 ;
    END
  END E1END[3]
  PIN E2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 96.600 225.000 97.200 ;
    END
  END E2BEG[0]
  PIN E2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 97.960 225.000 98.560 ;
    END
  END E2BEG[1]
  PIN E2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 99.320 225.000 99.920 ;
    END
  END E2BEG[2]
  PIN E2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 100.680 225.000 101.280 ;
    END
  END E2BEG[3]
  PIN E2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 102.040 225.000 102.640 ;
    END
  END E2BEG[4]
  PIN E2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 103.400 225.000 104.000 ;
    END
  END E2BEG[5]
  PIN E2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 104.760 225.000 105.360 ;
    END
  END E2BEG[6]
  PIN E2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 106.120 225.000 106.720 ;
    END
  END E2BEG[7]
  PIN E2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 107.480 225.000 108.080 ;
    END
  END E2BEGb[0]
  PIN E2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 108.840 225.000 109.440 ;
    END
  END E2BEGb[1]
  PIN E2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 110.200 225.000 110.800 ;
    END
  END E2BEGb[2]
  PIN E2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 111.560 225.000 112.160 ;
    END
  END E2BEGb[3]
  PIN E2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 112.920 225.000 113.520 ;
    END
  END E2BEGb[4]
  PIN E2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 114.280 225.000 114.880 ;
    END
  END E2BEGb[5]
  PIN E2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 115.640 225.000 116.240 ;
    END
  END E2BEGb[6]
  PIN E2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 117.000 225.000 117.600 ;
    END
  END E2BEGb[7]
  PIN E2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 0.800 108.080 ;
    END
  END E2END[0]
  PIN E2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 0.800 109.440 ;
    END
  END E2END[1]
  PIN E2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 0.800 110.800 ;
    END
  END E2END[2]
  PIN E2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.560 0.800 112.160 ;
    END
  END E2END[3]
  PIN E2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 0.800 113.520 ;
    END
  END E2END[4]
  PIN E2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.280 0.800 114.880 ;
    END
  END E2END[5]
  PIN E2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 0.800 116.240 ;
    END
  END E2END[6]
  PIN E2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 0.800 117.600 ;
    END
  END E2END[7]
  PIN E2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 0.800 97.200 ;
    END
  END E2MID[0]
  PIN E2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 0.800 98.560 ;
    END
  END E2MID[1]
  PIN E2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.320 0.800 99.920 ;
    END
  END E2MID[2]
  PIN E2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 0.800 101.280 ;
    END
  END E2MID[3]
  PIN E2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 0.800 102.640 ;
    END
  END E2MID[4]
  PIN E2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 0.800 104.000 ;
    END
  END E2MID[5]
  PIN E2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.760 0.800 105.360 ;
    END
  END E2MID[6]
  PIN E2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.120 0.800 106.720 ;
    END
  END E2MID[7]
  PIN E6BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 140.120 225.000 140.720 ;
    END
  END E6BEG[0]
  PIN E6BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 153.720 225.000 154.320 ;
    END
  END E6BEG[10]
  PIN E6BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 155.080 225.000 155.680 ;
    END
  END E6BEG[11]
  PIN E6BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 141.480 225.000 142.080 ;
    END
  END E6BEG[1]
  PIN E6BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 142.840 225.000 143.440 ;
    END
  END E6BEG[2]
  PIN E6BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 144.200 225.000 144.800 ;
    END
  END E6BEG[3]
  PIN E6BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 145.560 225.000 146.160 ;
    END
  END E6BEG[4]
  PIN E6BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 146.920 225.000 147.520 ;
    END
  END E6BEG[5]
  PIN E6BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 148.280 225.000 148.880 ;
    END
  END E6BEG[6]
  PIN E6BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 149.640 225.000 150.240 ;
    END
  END E6BEG[7]
  PIN E6BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 151.000 225.000 151.600 ;
    END
  END E6BEG[8]
  PIN E6BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 152.360 225.000 152.960 ;
    END
  END E6BEG[9]
  PIN E6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.120 0.800 140.720 ;
    END
  END E6END[0]
  PIN E6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.720 0.800 154.320 ;
    END
  END E6END[10]
  PIN E6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.080 0.800 155.680 ;
    END
  END E6END[11]
  PIN E6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.480 0.800 142.080 ;
    END
  END E6END[1]
  PIN E6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 0.800 143.440 ;
    END
  END E6END[2]
  PIN E6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.200 0.800 144.800 ;
    END
  END E6END[3]
  PIN E6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 0.800 146.160 ;
    END
  END E6END[4]
  PIN E6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.920 0.800 147.520 ;
    END
  END E6END[5]
  PIN E6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.280 0.800 148.880 ;
    END
  END E6END[6]
  PIN E6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 0.800 150.240 ;
    END
  END E6END[7]
  PIN E6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.000 0.800 151.600 ;
    END
  END E6END[8]
  PIN E6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.360 0.800 152.960 ;
    END
  END E6END[9]
  PIN EE4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 118.360 225.000 118.960 ;
    END
  END EE4BEG[0]
  PIN EE4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 131.960 225.000 132.560 ;
    END
  END EE4BEG[10]
  PIN EE4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 133.320 225.000 133.920 ;
    END
  END EE4BEG[11]
  PIN EE4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 134.680 225.000 135.280 ;
    END
  END EE4BEG[12]
  PIN EE4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 136.040 225.000 136.640 ;
    END
  END EE4BEG[13]
  PIN EE4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 137.400 225.000 138.000 ;
    END
  END EE4BEG[14]
  PIN EE4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 138.760 225.000 139.360 ;
    END
  END EE4BEG[15]
  PIN EE4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 119.720 225.000 120.320 ;
    END
  END EE4BEG[1]
  PIN EE4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 121.080 225.000 121.680 ;
    END
  END EE4BEG[2]
  PIN EE4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 122.440 225.000 123.040 ;
    END
  END EE4BEG[3]
  PIN EE4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 123.800 225.000 124.400 ;
    END
  END EE4BEG[4]
  PIN EE4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 125.160 225.000 125.760 ;
    END
  END EE4BEG[5]
  PIN EE4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 126.520 225.000 127.120 ;
    END
  END EE4BEG[6]
  PIN EE4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 127.880 225.000 128.480 ;
    END
  END EE4BEG[7]
  PIN EE4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 129.240 225.000 129.840 ;
    END
  END EE4BEG[8]
  PIN EE4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 130.600 225.000 131.200 ;
    END
  END EE4BEG[9]
  PIN EE4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.360 0.800 118.960 ;
    END
  END EE4END[0]
  PIN EE4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.960 0.800 132.560 ;
    END
  END EE4END[10]
  PIN EE4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.320 0.800 133.920 ;
    END
  END EE4END[11]
  PIN EE4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.680 0.800 135.280 ;
    END
  END EE4END[12]
  PIN EE4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 0.800 136.640 ;
    END
  END EE4END[13]
  PIN EE4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 0.800 138.000 ;
    END
  END EE4END[14]
  PIN EE4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.760 0.800 139.360 ;
    END
  END EE4END[15]
  PIN EE4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 0.800 120.320 ;
    END
  END EE4END[1]
  PIN EE4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 0.800 121.680 ;
    END
  END EE4END[2]
  PIN EE4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 0.800 123.040 ;
    END
  END EE4END[3]
  PIN EE4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.800 0.800 124.400 ;
    END
  END EE4END[4]
  PIN EE4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.160 0.800 125.760 ;
    END
  END EE4END[5]
  PIN EE4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 0.800 127.120 ;
    END
  END EE4END[6]
  PIN EE4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 0.800 128.480 ;
    END
  END EE4END[7]
  PIN EE4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 0.800 129.840 ;
    END
  END EE4END[8]
  PIN EE4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 0.800 131.200 ;
    END
  END EE4END[9]
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 0.800 157.040 ;
    END
  END FrameData[0]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 0.800 170.640 ;
    END
  END FrameData[10]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 171.400 0.800 172.000 ;
    END
  END FrameData[11]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.760 0.800 173.360 ;
    END
  END FrameData[12]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.120 0.800 174.720 ;
    END
  END FrameData[13]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.480 0.800 176.080 ;
    END
  END FrameData[14]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 0.800 177.440 ;
    END
  END FrameData[15]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.200 0.800 178.800 ;
    END
  END FrameData[16]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.560 0.800 180.160 ;
    END
  END FrameData[17]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.920 0.800 181.520 ;
    END
  END FrameData[18]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.280 0.800 182.880 ;
    END
  END FrameData[19]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.800 0.800 158.400 ;
    END
  END FrameData[1]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 0.800 184.240 ;
    END
  END FrameData[20]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.000 0.800 185.600 ;
    END
  END FrameData[21]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 186.360 0.800 186.960 ;
    END
  END FrameData[22]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.720 0.800 188.320 ;
    END
  END FrameData[23]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.080 0.800 189.680 ;
    END
  END FrameData[24]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 0.800 191.040 ;
    END
  END FrameData[25]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.800 0.800 192.400 ;
    END
  END FrameData[26]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 0.800 193.760 ;
    END
  END FrameData[27]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 194.520 0.800 195.120 ;
    END
  END FrameData[28]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.880 0.800 196.480 ;
    END
  END FrameData[29]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.160 0.800 159.760 ;
    END
  END FrameData[2]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 0.800 197.840 ;
    END
  END FrameData[30]
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.600 0.800 199.200 ;
    END
  END FrameData[31]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.520 0.800 161.120 ;
    END
  END FrameData[3]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.880 0.800 162.480 ;
    END
  END FrameData[4]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 0.800 163.840 ;
    END
  END FrameData[5]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.600 0.800 165.200 ;
    END
  END FrameData[6]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.960 0.800 166.560 ;
    END
  END FrameData[7]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 167.320 0.800 167.920 ;
    END
  END FrameData[8]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.680 0.800 169.280 ;
    END
  END FrameData[9]
  PIN FrameData_O[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 156.440 225.000 157.040 ;
    END
  END FrameData_O[0]
  PIN FrameData_O[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 170.040 225.000 170.640 ;
    END
  END FrameData_O[10]
  PIN FrameData_O[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 171.400 225.000 172.000 ;
    END
  END FrameData_O[11]
  PIN FrameData_O[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 172.760 225.000 173.360 ;
    END
  END FrameData_O[12]
  PIN FrameData_O[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 174.120 225.000 174.720 ;
    END
  END FrameData_O[13]
  PIN FrameData_O[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 175.480 225.000 176.080 ;
    END
  END FrameData_O[14]
  PIN FrameData_O[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 176.840 225.000 177.440 ;
    END
  END FrameData_O[15]
  PIN FrameData_O[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 178.200 225.000 178.800 ;
    END
  END FrameData_O[16]
  PIN FrameData_O[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 179.560 225.000 180.160 ;
    END
  END FrameData_O[17]
  PIN FrameData_O[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 180.920 225.000 181.520 ;
    END
  END FrameData_O[18]
  PIN FrameData_O[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 182.280 225.000 182.880 ;
    END
  END FrameData_O[19]
  PIN FrameData_O[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 157.800 225.000 158.400 ;
    END
  END FrameData_O[1]
  PIN FrameData_O[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 183.640 225.000 184.240 ;
    END
  END FrameData_O[20]
  PIN FrameData_O[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 185.000 225.000 185.600 ;
    END
  END FrameData_O[21]
  PIN FrameData_O[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 186.360 225.000 186.960 ;
    END
  END FrameData_O[22]
  PIN FrameData_O[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 187.720 225.000 188.320 ;
    END
  END FrameData_O[23]
  PIN FrameData_O[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 189.080 225.000 189.680 ;
    END
  END FrameData_O[24]
  PIN FrameData_O[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 190.440 225.000 191.040 ;
    END
  END FrameData_O[25]
  PIN FrameData_O[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 191.800 225.000 192.400 ;
    END
  END FrameData_O[26]
  PIN FrameData_O[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 193.160 225.000 193.760 ;
    END
  END FrameData_O[27]
  PIN FrameData_O[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 194.520 225.000 195.120 ;
    END
  END FrameData_O[28]
  PIN FrameData_O[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 195.880 225.000 196.480 ;
    END
  END FrameData_O[29]
  PIN FrameData_O[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 159.160 225.000 159.760 ;
    END
  END FrameData_O[2]
  PIN FrameData_O[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 197.240 225.000 197.840 ;
    END
  END FrameData_O[30]
  PIN FrameData_O[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 198.600 225.000 199.200 ;
    END
  END FrameData_O[31]
  PIN FrameData_O[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 160.520 225.000 161.120 ;
    END
  END FrameData_O[3]
  PIN FrameData_O[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 161.880 225.000 162.480 ;
    END
  END FrameData_O[4]
  PIN FrameData_O[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 163.240 225.000 163.840 ;
    END
  END FrameData_O[5]
  PIN FrameData_O[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 164.600 225.000 165.200 ;
    END
  END FrameData_O[6]
  PIN FrameData_O[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 165.960 225.000 166.560 ;
    END
  END FrameData_O[7]
  PIN FrameData_O[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 167.320 225.000 167.920 ;
    END
  END FrameData_O[8]
  PIN FrameData_O[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 168.680 225.000 169.280 ;
    END
  END FrameData_O[9]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 172.130 0.000 172.410 0.800 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 185.930 0.000 186.210 0.800 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 187.310 0.000 187.590 0.800 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 188.690 0.000 188.970 0.800 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 190.070 0.000 190.350 0.800 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 191.450 0.000 191.730 0.800 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 192.830 0.000 193.110 0.800 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 194.210 0.000 194.490 0.800 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 195.590 0.000 195.870 0.800 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 196.970 0.000 197.250 0.800 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 198.350 0.000 198.630 0.800 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 173.510 0.000 173.790 0.800 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 174.890 0.000 175.170 0.800 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 176.270 0.000 176.550 0.800 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 177.650 0.000 177.930 0.800 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 179.030 0.000 179.310 0.800 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 0.800 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 181.790 0.000 182.070 0.800 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 183.170 0.000 183.450 0.800 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 184.550 0.000 184.830 0.800 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 172.130 224.200 172.410 225.000 ;
    END
  END FrameStrobe_O[0]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 185.930 224.200 186.210 225.000 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 187.310 224.200 187.590 225.000 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 188.690 224.200 188.970 225.000 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 190.070 224.200 190.350 225.000 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 191.450 224.200 191.730 225.000 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 192.830 224.200 193.110 225.000 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 194.210 224.200 194.490 225.000 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 195.590 224.200 195.870 225.000 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 196.970 224.200 197.250 225.000 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 198.350 224.200 198.630 225.000 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 173.510 224.200 173.790 225.000 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 174.890 224.200 175.170 225.000 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 176.270 224.200 176.550 225.000 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 177.650 224.200 177.930 225.000 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 179.030 224.200 179.310 225.000 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 180.410 224.200 180.690 225.000 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 181.790 224.200 182.070 225.000 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 183.170 224.200 183.450 225.000 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 184.550 224.200 184.830 225.000 ;
    END
  END FrameStrobe_O[9]
  PIN N1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 25.850 224.200 26.130 225.000 ;
    END
  END N1BEG[0]
  PIN N1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 27.230 224.200 27.510 225.000 ;
    END
  END N1BEG[1]
  PIN N1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 28.610 224.200 28.890 225.000 ;
    END
  END N1BEG[2]
  PIN N1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 29.990 224.200 30.270 225.000 ;
    END
  END N1BEG[3]
  PIN N1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 0.800 ;
    END
  END N1END[0]
  PIN N1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 27.230 0.000 27.510 0.800 ;
    END
  END N1END[1]
  PIN N1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 28.610 0.000 28.890 0.800 ;
    END
  END N1END[2]
  PIN N1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 29.990 0.000 30.270 0.800 ;
    END
  END N1END[3]
  PIN N2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 31.370 224.200 31.650 225.000 ;
    END
  END N2BEG[0]
  PIN N2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 32.750 224.200 33.030 225.000 ;
    END
  END N2BEG[1]
  PIN N2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 34.130 224.200 34.410 225.000 ;
    END
  END N2BEG[2]
  PIN N2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 35.510 224.200 35.790 225.000 ;
    END
  END N2BEG[3]
  PIN N2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 36.890 224.200 37.170 225.000 ;
    END
  END N2BEG[4]
  PIN N2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 38.270 224.200 38.550 225.000 ;
    END
  END N2BEG[5]
  PIN N2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 39.650 224.200 39.930 225.000 ;
    END
  END N2BEG[6]
  PIN N2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 41.030 224.200 41.310 225.000 ;
    END
  END N2BEG[7]
  PIN N2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 42.410 224.200 42.690 225.000 ;
    END
  END N2BEGb[0]
  PIN N2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 43.790 224.200 44.070 225.000 ;
    END
  END N2BEGb[1]
  PIN N2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 45.170 224.200 45.450 225.000 ;
    END
  END N2BEGb[2]
  PIN N2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 46.550 224.200 46.830 225.000 ;
    END
  END N2BEGb[3]
  PIN N2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 47.930 224.200 48.210 225.000 ;
    END
  END N2BEGb[4]
  PIN N2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 49.310 224.200 49.590 225.000 ;
    END
  END N2BEGb[5]
  PIN N2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 50.690 224.200 50.970 225.000 ;
    END
  END N2BEGb[6]
  PIN N2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 52.070 224.200 52.350 225.000 ;
    END
  END N2BEGb[7]
  PIN N2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 42.410 0.000 42.690 0.800 ;
    END
  END N2END[0]
  PIN N2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 43.790 0.000 44.070 0.800 ;
    END
  END N2END[1]
  PIN N2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 0.800 ;
    END
  END N2END[2]
  PIN N2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 46.550 0.000 46.830 0.800 ;
    END
  END N2END[3]
  PIN N2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 47.930 0.000 48.210 0.800 ;
    END
  END N2END[4]
  PIN N2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 49.310 0.000 49.590 0.800 ;
    END
  END N2END[5]
  PIN N2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 50.690 0.000 50.970 0.800 ;
    END
  END N2END[6]
  PIN N2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 52.070 0.000 52.350 0.800 ;
    END
  END N2END[7]
  PIN N2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 31.370 0.000 31.650 0.800 ;
    END
  END N2MID[0]
  PIN N2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 32.750 0.000 33.030 0.800 ;
    END
  END N2MID[1]
  PIN N2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 34.130 0.000 34.410 0.800 ;
    END
  END N2MID[2]
  PIN N2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 0.800 ;
    END
  END N2MID[3]
  PIN N2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 36.890 0.000 37.170 0.800 ;
    END
  END N2MID[4]
  PIN N2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 38.270 0.000 38.550 0.800 ;
    END
  END N2MID[5]
  PIN N2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 39.650 0.000 39.930 0.800 ;
    END
  END N2MID[6]
  PIN N2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 41.030 0.000 41.310 0.800 ;
    END
  END N2MID[7]
  PIN N4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 53.450 224.200 53.730 225.000 ;
    END
  END N4BEG[0]
  PIN N4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 67.250 224.200 67.530 225.000 ;
    END
  END N4BEG[10]
  PIN N4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 68.630 224.200 68.910 225.000 ;
    END
  END N4BEG[11]
  PIN N4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 70.010 224.200 70.290 225.000 ;
    END
  END N4BEG[12]
  PIN N4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 71.390 224.200 71.670 225.000 ;
    END
  END N4BEG[13]
  PIN N4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 72.770 224.200 73.050 225.000 ;
    END
  END N4BEG[14]
  PIN N4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 74.150 224.200 74.430 225.000 ;
    END
  END N4BEG[15]
  PIN N4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 54.830 224.200 55.110 225.000 ;
    END
  END N4BEG[1]
  PIN N4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 56.210 224.200 56.490 225.000 ;
    END
  END N4BEG[2]
  PIN N4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 57.590 224.200 57.870 225.000 ;
    END
  END N4BEG[3]
  PIN N4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 58.970 224.200 59.250 225.000 ;
    END
  END N4BEG[4]
  PIN N4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 60.350 224.200 60.630 225.000 ;
    END
  END N4BEG[5]
  PIN N4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 61.730 224.200 62.010 225.000 ;
    END
  END N4BEG[6]
  PIN N4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 63.110 224.200 63.390 225.000 ;
    END
  END N4BEG[7]
  PIN N4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 64.490 224.200 64.770 225.000 ;
    END
  END N4BEG[8]
  PIN N4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 65.870 224.200 66.150 225.000 ;
    END
  END N4BEG[9]
  PIN N4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 53.450 0.000 53.730 0.800 ;
    END
  END N4END[0]
  PIN N4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 67.250 0.000 67.530 0.800 ;
    END
  END N4END[10]
  PIN N4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 68.630 0.000 68.910 0.800 ;
    END
  END N4END[11]
  PIN N4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 70.010 0.000 70.290 0.800 ;
    END
  END N4END[12]
  PIN N4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 71.390 0.000 71.670 0.800 ;
    END
  END N4END[13]
  PIN N4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 72.770 0.000 73.050 0.800 ;
    END
  END N4END[14]
  PIN N4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 0.800 ;
    END
  END N4END[15]
  PIN N4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 0.800 ;
    END
  END N4END[1]
  PIN N4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 56.210 0.000 56.490 0.800 ;
    END
  END N4END[2]
  PIN N4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 57.590 0.000 57.870 0.800 ;
    END
  END N4END[3]
  PIN N4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 58.970 0.000 59.250 0.800 ;
    END
  END N4END[4]
  PIN N4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 60.350 0.000 60.630 0.800 ;
    END
  END N4END[5]
  PIN N4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 61.730 0.000 62.010 0.800 ;
    END
  END N4END[6]
  PIN N4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 63.110 0.000 63.390 0.800 ;
    END
  END N4END[7]
  PIN N4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 0.800 ;
    END
  END N4END[8]
  PIN N4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 65.870 0.000 66.150 0.800 ;
    END
  END N4END[9]
  PIN NN4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 75.530 224.200 75.810 225.000 ;
    END
  END NN4BEG[0]
  PIN NN4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 89.330 224.200 89.610 225.000 ;
    END
  END NN4BEG[10]
  PIN NN4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 90.710 224.200 90.990 225.000 ;
    END
  END NN4BEG[11]
  PIN NN4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 92.090 224.200 92.370 225.000 ;
    END
  END NN4BEG[12]
  PIN NN4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 93.470 224.200 93.750 225.000 ;
    END
  END NN4BEG[13]
  PIN NN4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 94.850 224.200 95.130 225.000 ;
    END
  END NN4BEG[14]
  PIN NN4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 96.230 224.200 96.510 225.000 ;
    END
  END NN4BEG[15]
  PIN NN4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 76.910 224.200 77.190 225.000 ;
    END
  END NN4BEG[1]
  PIN NN4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 78.290 224.200 78.570 225.000 ;
    END
  END NN4BEG[2]
  PIN NN4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 79.670 224.200 79.950 225.000 ;
    END
  END NN4BEG[3]
  PIN NN4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 81.050 224.200 81.330 225.000 ;
    END
  END NN4BEG[4]
  PIN NN4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 82.430 224.200 82.710 225.000 ;
    END
  END NN4BEG[5]
  PIN NN4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 83.810 224.200 84.090 225.000 ;
    END
  END NN4BEG[6]
  PIN NN4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 85.190 224.200 85.470 225.000 ;
    END
  END NN4BEG[7]
  PIN NN4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 86.570 224.200 86.850 225.000 ;
    END
  END NN4BEG[8]
  PIN NN4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 87.950 224.200 88.230 225.000 ;
    END
  END NN4BEG[9]
  PIN NN4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 75.530 0.000 75.810 0.800 ;
    END
  END NN4END[0]
  PIN NN4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 89.330 0.000 89.610 0.800 ;
    END
  END NN4END[10]
  PIN NN4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 90.710 0.000 90.990 0.800 ;
    END
  END NN4END[11]
  PIN NN4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 92.090 0.000 92.370 0.800 ;
    END
  END NN4END[12]
  PIN NN4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 0.800 ;
    END
  END NN4END[13]
  PIN NN4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 94.850 0.000 95.130 0.800 ;
    END
  END NN4END[14]
  PIN NN4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 96.230 0.000 96.510 0.800 ;
    END
  END NN4END[15]
  PIN NN4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 76.910 0.000 77.190 0.800 ;
    END
  END NN4END[1]
  PIN NN4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 78.290 0.000 78.570 0.800 ;
    END
  END NN4END[2]
  PIN NN4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 79.670 0.000 79.950 0.800 ;
    END
  END NN4END[3]
  PIN NN4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 81.050 0.000 81.330 0.800 ;
    END
  END NN4END[4]
  PIN NN4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 82.430 0.000 82.710 0.800 ;
    END
  END NN4END[5]
  PIN NN4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 0.800 ;
    END
  END NN4END[6]
  PIN NN4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 85.190 0.000 85.470 0.800 ;
    END
  END NN4END[7]
  PIN NN4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 86.570 0.000 86.850 0.800 ;
    END
  END NN4END[8]
  PIN NN4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 87.950 0.000 88.230 0.800 ;
    END
  END NN4END[9]
  PIN S1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 97.610 0.000 97.890 0.800 ;
    END
  END S1BEG[0]
  PIN S1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 98.990 0.000 99.270 0.800 ;
    END
  END S1BEG[1]
  PIN S1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 100.370 0.000 100.650 0.800 ;
    END
  END S1BEG[2]
  PIN S1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 101.750 0.000 102.030 0.800 ;
    END
  END S1BEG[3]
  PIN S1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 97.610 224.200 97.890 225.000 ;
    END
  END S1END[0]
  PIN S1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 98.990 224.200 99.270 225.000 ;
    END
  END S1END[1]
  PIN S1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 100.370 224.200 100.650 225.000 ;
    END
  END S1END[2]
  PIN S1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 101.750 224.200 102.030 225.000 ;
    END
  END S1END[3]
  PIN S2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 114.170 0.000 114.450 0.800 ;
    END
  END S2BEG[0]
  PIN S2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 115.550 0.000 115.830 0.800 ;
    END
  END S2BEG[1]
  PIN S2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 116.930 0.000 117.210 0.800 ;
    END
  END S2BEG[2]
  PIN S2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 118.310 0.000 118.590 0.800 ;
    END
  END S2BEG[3]
  PIN S2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 0.800 ;
    END
  END S2BEG[4]
  PIN S2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 121.070 0.000 121.350 0.800 ;
    END
  END S2BEG[5]
  PIN S2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 0.800 ;
    END
  END S2BEG[6]
  PIN S2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 123.830 0.000 124.110 0.800 ;
    END
  END S2BEG[7]
  PIN S2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 0.800 ;
    END
  END S2BEGb[0]
  PIN S2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 104.510 0.000 104.790 0.800 ;
    END
  END S2BEGb[1]
  PIN S2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 105.890 0.000 106.170 0.800 ;
    END
  END S2BEGb[2]
  PIN S2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 107.270 0.000 107.550 0.800 ;
    END
  END S2BEGb[3]
  PIN S2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 108.650 0.000 108.930 0.800 ;
    END
  END S2BEGb[4]
  PIN S2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 110.030 0.000 110.310 0.800 ;
    END
  END S2BEGb[5]
  PIN S2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 111.410 0.000 111.690 0.800 ;
    END
  END S2BEGb[6]
  PIN S2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 0.800 ;
    END
  END S2BEGb[7]
  PIN S2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 103.130 224.200 103.410 225.000 ;
    END
  END S2END[0]
  PIN S2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 104.510 224.200 104.790 225.000 ;
    END
  END S2END[1]
  PIN S2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 105.890 224.200 106.170 225.000 ;
    END
  END S2END[2]
  PIN S2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 107.270 224.200 107.550 225.000 ;
    END
  END S2END[3]
  PIN S2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 108.650 224.200 108.930 225.000 ;
    END
  END S2END[4]
  PIN S2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 110.030 224.200 110.310 225.000 ;
    END
  END S2END[5]
  PIN S2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 111.410 224.200 111.690 225.000 ;
    END
  END S2END[6]
  PIN S2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 112.790 224.200 113.070 225.000 ;
    END
  END S2END[7]
  PIN S2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 114.170 224.200 114.450 225.000 ;
    END
  END S2MID[0]
  PIN S2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 115.550 224.200 115.830 225.000 ;
    END
  END S2MID[1]
  PIN S2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 116.930 224.200 117.210 225.000 ;
    END
  END S2MID[2]
  PIN S2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 118.310 224.200 118.590 225.000 ;
    END
  END S2MID[3]
  PIN S2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 119.690 224.200 119.970 225.000 ;
    END
  END S2MID[4]
  PIN S2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 121.070 224.200 121.350 225.000 ;
    END
  END S2MID[5]
  PIN S2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 122.450 224.200 122.730 225.000 ;
    END
  END S2MID[6]
  PIN S2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 123.830 224.200 124.110 225.000 ;
    END
  END S2MID[7]
  PIN S4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 125.210 0.000 125.490 0.800 ;
    END
  END S4BEG[0]
  PIN S4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 139.010 0.000 139.290 0.800 ;
    END
  END S4BEG[10]
  PIN S4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 140.390 0.000 140.670 0.800 ;
    END
  END S4BEG[11]
  PIN S4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 0.800 ;
    END
  END S4BEG[12]
  PIN S4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 143.150 0.000 143.430 0.800 ;
    END
  END S4BEG[13]
  PIN S4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 144.530 0.000 144.810 0.800 ;
    END
  END S4BEG[14]
  PIN S4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 145.910 0.000 146.190 0.800 ;
    END
  END S4BEG[15]
  PIN S4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 126.590 0.000 126.870 0.800 ;
    END
  END S4BEG[1]
  PIN S4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 127.970 0.000 128.250 0.800 ;
    END
  END S4BEG[2]
  PIN S4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 129.350 0.000 129.630 0.800 ;
    END
  END S4BEG[3]
  PIN S4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 130.730 0.000 131.010 0.800 ;
    END
  END S4BEG[4]
  PIN S4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 0.800 ;
    END
  END S4BEG[5]
  PIN S4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 133.490 0.000 133.770 0.800 ;
    END
  END S4BEG[6]
  PIN S4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 134.870 0.000 135.150 0.800 ;
    END
  END S4BEG[7]
  PIN S4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 136.250 0.000 136.530 0.800 ;
    END
  END S4BEG[8]
  PIN S4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 137.630 0.000 137.910 0.800 ;
    END
  END S4BEG[9]
  PIN S4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 125.210 224.200 125.490 225.000 ;
    END
  END S4END[0]
  PIN S4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 139.010 224.200 139.290 225.000 ;
    END
  END S4END[10]
  PIN S4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 140.390 224.200 140.670 225.000 ;
    END
  END S4END[11]
  PIN S4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 141.770 224.200 142.050 225.000 ;
    END
  END S4END[12]
  PIN S4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 143.150 224.200 143.430 225.000 ;
    END
  END S4END[13]
  PIN S4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 144.530 224.200 144.810 225.000 ;
    END
  END S4END[14]
  PIN S4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 145.910 224.200 146.190 225.000 ;
    END
  END S4END[15]
  PIN S4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 126.590 224.200 126.870 225.000 ;
    END
  END S4END[1]
  PIN S4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 127.970 224.200 128.250 225.000 ;
    END
  END S4END[2]
  PIN S4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 129.350 224.200 129.630 225.000 ;
    END
  END S4END[3]
  PIN S4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 130.730 224.200 131.010 225.000 ;
    END
  END S4END[4]
  PIN S4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 132.110 224.200 132.390 225.000 ;
    END
  END S4END[5]
  PIN S4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 133.490 224.200 133.770 225.000 ;
    END
  END S4END[6]
  PIN S4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 134.870 224.200 135.150 225.000 ;
    END
  END S4END[7]
  PIN S4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 136.250 224.200 136.530 225.000 ;
    END
  END S4END[8]
  PIN S4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 137.630 224.200 137.910 225.000 ;
    END
  END S4END[9]
  PIN SS4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 147.290 0.000 147.570 0.800 ;
    END
  END SS4BEG[0]
  PIN SS4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 0.800 ;
    END
  END SS4BEG[10]
  PIN SS4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 162.470 0.000 162.750 0.800 ;
    END
  END SS4BEG[11]
  PIN SS4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 163.850 0.000 164.130 0.800 ;
    END
  END SS4BEG[12]
  PIN SS4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 165.230 0.000 165.510 0.800 ;
    END
  END SS4BEG[13]
  PIN SS4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 166.610 0.000 166.890 0.800 ;
    END
  END SS4BEG[14]
  PIN SS4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 167.990 0.000 168.270 0.800 ;
    END
  END SS4BEG[15]
  PIN SS4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 148.670 0.000 148.950 0.800 ;
    END
  END SS4BEG[1]
  PIN SS4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 150.050 0.000 150.330 0.800 ;
    END
  END SS4BEG[2]
  PIN SS4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 151.430 0.000 151.710 0.800 ;
    END
  END SS4BEG[3]
  PIN SS4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 152.810 0.000 153.090 0.800 ;
    END
  END SS4BEG[4]
  PIN SS4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 154.190 0.000 154.470 0.800 ;
    END
  END SS4BEG[5]
  PIN SS4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 155.570 0.000 155.850 0.800 ;
    END
  END SS4BEG[6]
  PIN SS4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 156.950 0.000 157.230 0.800 ;
    END
  END SS4BEG[7]
  PIN SS4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 158.330 0.000 158.610 0.800 ;
    END
  END SS4BEG[8]
  PIN SS4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 159.710 0.000 159.990 0.800 ;
    END
  END SS4BEG[9]
  PIN SS4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 147.290 224.200 147.570 225.000 ;
    END
  END SS4END[0]
  PIN SS4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 161.090 224.200 161.370 225.000 ;
    END
  END SS4END[10]
  PIN SS4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 162.470 224.200 162.750 225.000 ;
    END
  END SS4END[11]
  PIN SS4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 163.850 224.200 164.130 225.000 ;
    END
  END SS4END[12]
  PIN SS4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 165.230 224.200 165.510 225.000 ;
    END
  END SS4END[13]
  PIN SS4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 166.610 224.200 166.890 225.000 ;
    END
  END SS4END[14]
  PIN SS4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 167.990 224.200 168.270 225.000 ;
    END
  END SS4END[15]
  PIN SS4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 148.670 224.200 148.950 225.000 ;
    END
  END SS4END[1]
  PIN SS4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 150.050 224.200 150.330 225.000 ;
    END
  END SS4END[2]
  PIN SS4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 151.430 224.200 151.710 225.000 ;
    END
  END SS4END[3]
  PIN SS4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 152.810 224.200 153.090 225.000 ;
    END
  END SS4END[4]
  PIN SS4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 154.190 224.200 154.470 225.000 ;
    END
  END SS4END[5]
  PIN SS4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 155.570 224.200 155.850 225.000 ;
    END
  END SS4END[6]
  PIN SS4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 156.950 224.200 157.230 225.000 ;
    END
  END SS4END[7]
  PIN SS4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 158.330 224.200 158.610 225.000 ;
    END
  END SS4END[8]
  PIN SS4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 159.710 224.200 159.990 225.000 ;
    END
  END SS4END[9]
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.124000 ;
    PORT
      LAYER met2 ;
        RECT 169.370 0.000 169.650 0.800 ;
    END
  END UserCLK
  PIN UserCLKo
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 169.370 224.200 169.650 225.000 ;
    END
  END UserCLKo
  PIN W1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 0.800 26.480 ;
    END
  END W1BEG[0]
  PIN W1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 0.800 27.840 ;
    END
  END W1BEG[1]
  PIN W1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 0.800 29.200 ;
    END
  END W1BEG[2]
  PIN W1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 0.800 30.560 ;
    END
  END W1BEG[3]
  PIN W1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 25.880 225.000 26.480 ;
    END
  END W1END[0]
  PIN W1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 27.240 225.000 27.840 ;
    END
  END W1END[1]
  PIN W1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 28.600 225.000 29.200 ;
    END
  END W1END[2]
  PIN W1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 29.960 225.000 30.560 ;
    END
  END W1END[3]
  PIN W2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 0.800 31.920 ;
    END
  END W2BEG[0]
  PIN W2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 0.800 33.280 ;
    END
  END W2BEG[1]
  PIN W2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 0.800 34.640 ;
    END
  END W2BEG[2]
  PIN W2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 0.800 36.000 ;
    END
  END W2BEG[3]
  PIN W2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.760 0.800 37.360 ;
    END
  END W2BEG[4]
  PIN W2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 0.800 38.720 ;
    END
  END W2BEG[5]
  PIN W2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 0.800 40.080 ;
    END
  END W2BEG[6]
  PIN W2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 0.800 41.440 ;
    END
  END W2BEG[7]
  PIN W2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 0.800 42.800 ;
    END
  END W2BEGb[0]
  PIN W2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 0.800 44.160 ;
    END
  END W2BEGb[1]
  PIN W2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 0.800 45.520 ;
    END
  END W2BEGb[2]
  PIN W2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 0.800 46.880 ;
    END
  END W2BEGb[3]
  PIN W2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 0.800 48.240 ;
    END
  END W2BEGb[4]
  PIN W2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 0.800 49.600 ;
    END
  END W2BEGb[5]
  PIN W2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 0.800 50.960 ;
    END
  END W2BEGb[6]
  PIN W2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 0.800 52.320 ;
    END
  END W2BEGb[7]
  PIN W2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 42.200 225.000 42.800 ;
    END
  END W2END[0]
  PIN W2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 43.560 225.000 44.160 ;
    END
  END W2END[1]
  PIN W2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 44.920 225.000 45.520 ;
    END
  END W2END[2]
  PIN W2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 46.280 225.000 46.880 ;
    END
  END W2END[3]
  PIN W2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 47.640 225.000 48.240 ;
    END
  END W2END[4]
  PIN W2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 49.000 225.000 49.600 ;
    END
  END W2END[5]
  PIN W2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 50.360 225.000 50.960 ;
    END
  END W2END[6]
  PIN W2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 51.720 225.000 52.320 ;
    END
  END W2END[7]
  PIN W2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 31.320 225.000 31.920 ;
    END
  END W2MID[0]
  PIN W2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 32.680 225.000 33.280 ;
    END
  END W2MID[1]
  PIN W2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 34.040 225.000 34.640 ;
    END
  END W2MID[2]
  PIN W2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 35.400 225.000 36.000 ;
    END
  END W2MID[3]
  PIN W2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 36.760 225.000 37.360 ;
    END
  END W2MID[4]
  PIN W2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 38.120 225.000 38.720 ;
    END
  END W2MID[5]
  PIN W2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 39.480 225.000 40.080 ;
    END
  END W2MID[6]
  PIN W2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 40.840 225.000 41.440 ;
    END
  END W2MID[7]
  PIN W6BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 0.800 75.440 ;
    END
  END W6BEG[0]
  PIN W6BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 0.800 89.040 ;
    END
  END W6BEG[10]
  PIN W6BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 0.800 90.400 ;
    END
  END W6BEG[11]
  PIN W6BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 0.800 76.800 ;
    END
  END W6BEG[1]
  PIN W6BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.560 0.800 78.160 ;
    END
  END W6BEG[2]
  PIN W6BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 0.800 79.520 ;
    END
  END W6BEG[3]
  PIN W6BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 0.800 80.880 ;
    END
  END W6BEG[4]
  PIN W6BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 0.800 82.240 ;
    END
  END W6BEG[5]
  PIN W6BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 0.800 83.600 ;
    END
  END W6BEG[6]
  PIN W6BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 0.800 84.960 ;
    END
  END W6BEG[7]
  PIN W6BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 0.800 86.320 ;
    END
  END W6BEG[8]
  PIN W6BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 0.800 87.680 ;
    END
  END W6BEG[9]
  PIN W6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 74.840 225.000 75.440 ;
    END
  END W6END[0]
  PIN W6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 88.440 225.000 89.040 ;
    END
  END W6END[10]
  PIN W6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 89.800 225.000 90.400 ;
    END
  END W6END[11]
  PIN W6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 76.200 225.000 76.800 ;
    END
  END W6END[1]
  PIN W6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 77.560 225.000 78.160 ;
    END
  END W6END[2]
  PIN W6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 78.920 225.000 79.520 ;
    END
  END W6END[3]
  PIN W6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 80.280 225.000 80.880 ;
    END
  END W6END[4]
  PIN W6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 81.640 225.000 82.240 ;
    END
  END W6END[5]
  PIN W6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 83.000 225.000 83.600 ;
    END
  END W6END[6]
  PIN W6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 84.360 225.000 84.960 ;
    END
  END W6END[7]
  PIN W6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 85.720 225.000 86.320 ;
    END
  END W6END[8]
  PIN W6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 87.080 225.000 87.680 ;
    END
  END W6END[9]
  PIN WW4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 0.800 53.680 ;
    END
  END WW4BEG[0]
  PIN WW4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.680 0.800 67.280 ;
    END
  END WW4BEG[10]
  PIN WW4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 0.800 68.640 ;
    END
  END WW4BEG[11]
  PIN WW4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 0.800 70.000 ;
    END
  END WW4BEG[12]
  PIN WW4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 0.800 71.360 ;
    END
  END WW4BEG[13]
  PIN WW4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 0.800 72.720 ;
    END
  END WW4BEG[14]
  PIN WW4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.480 0.800 74.080 ;
    END
  END WW4BEG[15]
  PIN WW4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 0.800 55.040 ;
    END
  END WW4BEG[1]
  PIN WW4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 0.800 56.400 ;
    END
  END WW4BEG[2]
  PIN WW4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 0.800 57.760 ;
    END
  END WW4BEG[3]
  PIN WW4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 0.800 59.120 ;
    END
  END WW4BEG[4]
  PIN WW4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 0.800 60.480 ;
    END
  END WW4BEG[5]
  PIN WW4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 0.800 61.840 ;
    END
  END WW4BEG[6]
  PIN WW4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 0.800 63.200 ;
    END
  END WW4BEG[7]
  PIN WW4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 0.800 64.560 ;
    END
  END WW4BEG[8]
  PIN WW4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 0.800 65.920 ;
    END
  END WW4BEG[9]
  PIN WW4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 53.080 225.000 53.680 ;
    END
  END WW4END[0]
  PIN WW4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 66.680 225.000 67.280 ;
    END
  END WW4END[10]
  PIN WW4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 68.040 225.000 68.640 ;
    END
  END WW4END[11]
  PIN WW4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 69.400 225.000 70.000 ;
    END
  END WW4END[12]
  PIN WW4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 70.760 225.000 71.360 ;
    END
  END WW4END[13]
  PIN WW4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 72.120 225.000 72.720 ;
    END
  END WW4END[14]
  PIN WW4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 73.480 225.000 74.080 ;
    END
  END WW4END[15]
  PIN WW4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 54.440 225.000 55.040 ;
    END
  END WW4END[1]
  PIN WW4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 55.800 225.000 56.400 ;
    END
  END WW4END[2]
  PIN WW4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 57.160 225.000 57.760 ;
    END
  END WW4END[3]
  PIN WW4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 58.520 225.000 59.120 ;
    END
  END WW4END[4]
  PIN WW4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 59.880 225.000 60.480 ;
    END
  END WW4END[5]
  PIN WW4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 61.240 225.000 61.840 ;
    END
  END WW4END[6]
  PIN WW4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 62.600 225.000 63.200 ;
    END
  END WW4END[7]
  PIN WW4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 63.960 225.000 64.560 ;
    END
  END WW4END[8]
  PIN WW4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 65.320 225.000 65.920 ;
    END
  END WW4END[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 17.820 5.200 19.420 217.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 92.820 5.200 94.420 217.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 167.820 5.200 169.420 217.840 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 55.320 5.200 56.920 217.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 130.320 5.200 131.920 217.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 205.320 5.200 206.920 217.840 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 2.300 5.355 222.640 217.685 ;
      LAYER met1 ;
        RECT 0.070 0.380 224.870 224.020 ;
      LAYER met2 ;
        RECT 0.100 223.920 25.570 224.810 ;
        RECT 26.410 223.920 26.950 224.810 ;
        RECT 27.790 223.920 28.330 224.810 ;
        RECT 29.170 223.920 29.710 224.810 ;
        RECT 30.550 223.920 31.090 224.810 ;
        RECT 31.930 223.920 32.470 224.810 ;
        RECT 33.310 223.920 33.850 224.810 ;
        RECT 34.690 223.920 35.230 224.810 ;
        RECT 36.070 223.920 36.610 224.810 ;
        RECT 37.450 223.920 37.990 224.810 ;
        RECT 38.830 223.920 39.370 224.810 ;
        RECT 40.210 223.920 40.750 224.810 ;
        RECT 41.590 223.920 42.130 224.810 ;
        RECT 42.970 223.920 43.510 224.810 ;
        RECT 44.350 223.920 44.890 224.810 ;
        RECT 45.730 223.920 46.270 224.810 ;
        RECT 47.110 223.920 47.650 224.810 ;
        RECT 48.490 223.920 49.030 224.810 ;
        RECT 49.870 223.920 50.410 224.810 ;
        RECT 51.250 223.920 51.790 224.810 ;
        RECT 52.630 223.920 53.170 224.810 ;
        RECT 54.010 223.920 54.550 224.810 ;
        RECT 55.390 223.920 55.930 224.810 ;
        RECT 56.770 223.920 57.310 224.810 ;
        RECT 58.150 223.920 58.690 224.810 ;
        RECT 59.530 223.920 60.070 224.810 ;
        RECT 60.910 223.920 61.450 224.810 ;
        RECT 62.290 223.920 62.830 224.810 ;
        RECT 63.670 223.920 64.210 224.810 ;
        RECT 65.050 223.920 65.590 224.810 ;
        RECT 66.430 223.920 66.970 224.810 ;
        RECT 67.810 223.920 68.350 224.810 ;
        RECT 69.190 223.920 69.730 224.810 ;
        RECT 70.570 223.920 71.110 224.810 ;
        RECT 71.950 223.920 72.490 224.810 ;
        RECT 73.330 223.920 73.870 224.810 ;
        RECT 74.710 223.920 75.250 224.810 ;
        RECT 76.090 223.920 76.630 224.810 ;
        RECT 77.470 223.920 78.010 224.810 ;
        RECT 78.850 223.920 79.390 224.810 ;
        RECT 80.230 223.920 80.770 224.810 ;
        RECT 81.610 223.920 82.150 224.810 ;
        RECT 82.990 223.920 83.530 224.810 ;
        RECT 84.370 223.920 84.910 224.810 ;
        RECT 85.750 223.920 86.290 224.810 ;
        RECT 87.130 223.920 87.670 224.810 ;
        RECT 88.510 223.920 89.050 224.810 ;
        RECT 89.890 223.920 90.430 224.810 ;
        RECT 91.270 223.920 91.810 224.810 ;
        RECT 92.650 223.920 93.190 224.810 ;
        RECT 94.030 223.920 94.570 224.810 ;
        RECT 95.410 223.920 95.950 224.810 ;
        RECT 96.790 223.920 97.330 224.810 ;
        RECT 98.170 223.920 98.710 224.810 ;
        RECT 99.550 223.920 100.090 224.810 ;
        RECT 100.930 223.920 101.470 224.810 ;
        RECT 102.310 223.920 102.850 224.810 ;
        RECT 103.690 223.920 104.230 224.810 ;
        RECT 105.070 223.920 105.610 224.810 ;
        RECT 106.450 223.920 106.990 224.810 ;
        RECT 107.830 223.920 108.370 224.810 ;
        RECT 109.210 223.920 109.750 224.810 ;
        RECT 110.590 223.920 111.130 224.810 ;
        RECT 111.970 223.920 112.510 224.810 ;
        RECT 113.350 223.920 113.890 224.810 ;
        RECT 114.730 223.920 115.270 224.810 ;
        RECT 116.110 223.920 116.650 224.810 ;
        RECT 117.490 223.920 118.030 224.810 ;
        RECT 118.870 223.920 119.410 224.810 ;
        RECT 120.250 223.920 120.790 224.810 ;
        RECT 121.630 223.920 122.170 224.810 ;
        RECT 123.010 223.920 123.550 224.810 ;
        RECT 124.390 223.920 124.930 224.810 ;
        RECT 125.770 223.920 126.310 224.810 ;
        RECT 127.150 223.920 127.690 224.810 ;
        RECT 128.530 223.920 129.070 224.810 ;
        RECT 129.910 223.920 130.450 224.810 ;
        RECT 131.290 223.920 131.830 224.810 ;
        RECT 132.670 223.920 133.210 224.810 ;
        RECT 134.050 223.920 134.590 224.810 ;
        RECT 135.430 223.920 135.970 224.810 ;
        RECT 136.810 223.920 137.350 224.810 ;
        RECT 138.190 223.920 138.730 224.810 ;
        RECT 139.570 223.920 140.110 224.810 ;
        RECT 140.950 223.920 141.490 224.810 ;
        RECT 142.330 223.920 142.870 224.810 ;
        RECT 143.710 223.920 144.250 224.810 ;
        RECT 145.090 223.920 145.630 224.810 ;
        RECT 146.470 223.920 147.010 224.810 ;
        RECT 147.850 223.920 148.390 224.810 ;
        RECT 149.230 223.920 149.770 224.810 ;
        RECT 150.610 223.920 151.150 224.810 ;
        RECT 151.990 223.920 152.530 224.810 ;
        RECT 153.370 223.920 153.910 224.810 ;
        RECT 154.750 223.920 155.290 224.810 ;
        RECT 156.130 223.920 156.670 224.810 ;
        RECT 157.510 223.920 158.050 224.810 ;
        RECT 158.890 223.920 159.430 224.810 ;
        RECT 160.270 223.920 160.810 224.810 ;
        RECT 161.650 223.920 162.190 224.810 ;
        RECT 163.030 223.920 163.570 224.810 ;
        RECT 164.410 223.920 164.950 224.810 ;
        RECT 165.790 223.920 166.330 224.810 ;
        RECT 167.170 223.920 167.710 224.810 ;
        RECT 168.550 223.920 169.090 224.810 ;
        RECT 169.930 223.920 170.470 224.810 ;
        RECT 171.310 223.920 171.850 224.810 ;
        RECT 172.690 223.920 173.230 224.810 ;
        RECT 174.070 223.920 174.610 224.810 ;
        RECT 175.450 223.920 175.990 224.810 ;
        RECT 176.830 223.920 177.370 224.810 ;
        RECT 178.210 223.920 178.750 224.810 ;
        RECT 179.590 223.920 180.130 224.810 ;
        RECT 180.970 223.920 181.510 224.810 ;
        RECT 182.350 223.920 182.890 224.810 ;
        RECT 183.730 223.920 184.270 224.810 ;
        RECT 185.110 223.920 185.650 224.810 ;
        RECT 186.490 223.920 187.030 224.810 ;
        RECT 187.870 223.920 188.410 224.810 ;
        RECT 189.250 223.920 189.790 224.810 ;
        RECT 190.630 223.920 191.170 224.810 ;
        RECT 192.010 223.920 192.550 224.810 ;
        RECT 193.390 223.920 193.930 224.810 ;
        RECT 194.770 223.920 195.310 224.810 ;
        RECT 196.150 223.920 196.690 224.810 ;
        RECT 197.530 223.920 198.070 224.810 ;
        RECT 198.910 223.920 224.850 224.810 ;
        RECT 0.100 1.080 224.850 223.920 ;
        RECT 0.100 0.270 25.570 1.080 ;
        RECT 26.410 0.270 26.950 1.080 ;
        RECT 27.790 0.270 28.330 1.080 ;
        RECT 29.170 0.270 29.710 1.080 ;
        RECT 30.550 0.270 31.090 1.080 ;
        RECT 31.930 0.270 32.470 1.080 ;
        RECT 33.310 0.270 33.850 1.080 ;
        RECT 34.690 0.270 35.230 1.080 ;
        RECT 36.070 0.270 36.610 1.080 ;
        RECT 37.450 0.270 37.990 1.080 ;
        RECT 38.830 0.270 39.370 1.080 ;
        RECT 40.210 0.270 40.750 1.080 ;
        RECT 41.590 0.270 42.130 1.080 ;
        RECT 42.970 0.270 43.510 1.080 ;
        RECT 44.350 0.270 44.890 1.080 ;
        RECT 45.730 0.270 46.270 1.080 ;
        RECT 47.110 0.270 47.650 1.080 ;
        RECT 48.490 0.270 49.030 1.080 ;
        RECT 49.870 0.270 50.410 1.080 ;
        RECT 51.250 0.270 51.790 1.080 ;
        RECT 52.630 0.270 53.170 1.080 ;
        RECT 54.010 0.270 54.550 1.080 ;
        RECT 55.390 0.270 55.930 1.080 ;
        RECT 56.770 0.270 57.310 1.080 ;
        RECT 58.150 0.270 58.690 1.080 ;
        RECT 59.530 0.270 60.070 1.080 ;
        RECT 60.910 0.270 61.450 1.080 ;
        RECT 62.290 0.270 62.830 1.080 ;
        RECT 63.670 0.270 64.210 1.080 ;
        RECT 65.050 0.270 65.590 1.080 ;
        RECT 66.430 0.270 66.970 1.080 ;
        RECT 67.810 0.270 68.350 1.080 ;
        RECT 69.190 0.270 69.730 1.080 ;
        RECT 70.570 0.270 71.110 1.080 ;
        RECT 71.950 0.270 72.490 1.080 ;
        RECT 73.330 0.270 73.870 1.080 ;
        RECT 74.710 0.270 75.250 1.080 ;
        RECT 76.090 0.270 76.630 1.080 ;
        RECT 77.470 0.270 78.010 1.080 ;
        RECT 78.850 0.270 79.390 1.080 ;
        RECT 80.230 0.270 80.770 1.080 ;
        RECT 81.610 0.270 82.150 1.080 ;
        RECT 82.990 0.270 83.530 1.080 ;
        RECT 84.370 0.270 84.910 1.080 ;
        RECT 85.750 0.270 86.290 1.080 ;
        RECT 87.130 0.270 87.670 1.080 ;
        RECT 88.510 0.270 89.050 1.080 ;
        RECT 89.890 0.270 90.430 1.080 ;
        RECT 91.270 0.270 91.810 1.080 ;
        RECT 92.650 0.270 93.190 1.080 ;
        RECT 94.030 0.270 94.570 1.080 ;
        RECT 95.410 0.270 95.950 1.080 ;
        RECT 96.790 0.270 97.330 1.080 ;
        RECT 98.170 0.270 98.710 1.080 ;
        RECT 99.550 0.270 100.090 1.080 ;
        RECT 100.930 0.270 101.470 1.080 ;
        RECT 102.310 0.270 102.850 1.080 ;
        RECT 103.690 0.270 104.230 1.080 ;
        RECT 105.070 0.270 105.610 1.080 ;
        RECT 106.450 0.270 106.990 1.080 ;
        RECT 107.830 0.270 108.370 1.080 ;
        RECT 109.210 0.270 109.750 1.080 ;
        RECT 110.590 0.270 111.130 1.080 ;
        RECT 111.970 0.270 112.510 1.080 ;
        RECT 113.350 0.270 113.890 1.080 ;
        RECT 114.730 0.270 115.270 1.080 ;
        RECT 116.110 0.270 116.650 1.080 ;
        RECT 117.490 0.270 118.030 1.080 ;
        RECT 118.870 0.270 119.410 1.080 ;
        RECT 120.250 0.270 120.790 1.080 ;
        RECT 121.630 0.270 122.170 1.080 ;
        RECT 123.010 0.270 123.550 1.080 ;
        RECT 124.390 0.270 124.930 1.080 ;
        RECT 125.770 0.270 126.310 1.080 ;
        RECT 127.150 0.270 127.690 1.080 ;
        RECT 128.530 0.270 129.070 1.080 ;
        RECT 129.910 0.270 130.450 1.080 ;
        RECT 131.290 0.270 131.830 1.080 ;
        RECT 132.670 0.270 133.210 1.080 ;
        RECT 134.050 0.270 134.590 1.080 ;
        RECT 135.430 0.270 135.970 1.080 ;
        RECT 136.810 0.270 137.350 1.080 ;
        RECT 138.190 0.270 138.730 1.080 ;
        RECT 139.570 0.270 140.110 1.080 ;
        RECT 140.950 0.270 141.490 1.080 ;
        RECT 142.330 0.270 142.870 1.080 ;
        RECT 143.710 0.270 144.250 1.080 ;
        RECT 145.090 0.270 145.630 1.080 ;
        RECT 146.470 0.270 147.010 1.080 ;
        RECT 147.850 0.270 148.390 1.080 ;
        RECT 149.230 0.270 149.770 1.080 ;
        RECT 150.610 0.270 151.150 1.080 ;
        RECT 151.990 0.270 152.530 1.080 ;
        RECT 153.370 0.270 153.910 1.080 ;
        RECT 154.750 0.270 155.290 1.080 ;
        RECT 156.130 0.270 156.670 1.080 ;
        RECT 157.510 0.270 158.050 1.080 ;
        RECT 158.890 0.270 159.430 1.080 ;
        RECT 160.270 0.270 160.810 1.080 ;
        RECT 161.650 0.270 162.190 1.080 ;
        RECT 163.030 0.270 163.570 1.080 ;
        RECT 164.410 0.270 164.950 1.080 ;
        RECT 165.790 0.270 166.330 1.080 ;
        RECT 167.170 0.270 167.710 1.080 ;
        RECT 168.550 0.270 169.090 1.080 ;
        RECT 169.930 0.270 170.470 1.080 ;
        RECT 171.310 0.270 171.850 1.080 ;
        RECT 172.690 0.270 173.230 1.080 ;
        RECT 174.070 0.270 174.610 1.080 ;
        RECT 175.450 0.270 175.990 1.080 ;
        RECT 176.830 0.270 177.370 1.080 ;
        RECT 178.210 0.270 178.750 1.080 ;
        RECT 179.590 0.270 180.130 1.080 ;
        RECT 180.970 0.270 181.510 1.080 ;
        RECT 182.350 0.270 182.890 1.080 ;
        RECT 183.730 0.270 184.270 1.080 ;
        RECT 185.110 0.270 185.650 1.080 ;
        RECT 186.490 0.270 187.030 1.080 ;
        RECT 187.870 0.270 188.410 1.080 ;
        RECT 189.250 0.270 189.790 1.080 ;
        RECT 190.630 0.270 191.170 1.080 ;
        RECT 192.010 0.270 192.550 1.080 ;
        RECT 193.390 0.270 193.930 1.080 ;
        RECT 194.770 0.270 195.310 1.080 ;
        RECT 196.150 0.270 196.690 1.080 ;
        RECT 197.530 0.270 198.070 1.080 ;
        RECT 198.910 0.270 224.850 1.080 ;
      LAYER met3 ;
        RECT 0.800 199.600 224.875 219.465 ;
        RECT 1.200 25.480 223.800 199.600 ;
        RECT 0.800 0.855 224.875 25.480 ;
      LAYER met4 ;
        RECT 1.215 218.240 223.265 219.465 ;
        RECT 1.215 4.800 17.420 218.240 ;
        RECT 19.820 4.800 54.920 218.240 ;
        RECT 57.320 4.800 92.420 218.240 ;
        RECT 94.820 4.800 129.920 218.240 ;
        RECT 132.320 4.800 167.420 218.240 ;
        RECT 169.820 4.800 204.920 218.240 ;
        RECT 207.320 4.800 223.265 218.240 ;
        RECT 1.215 1.535 223.265 4.800 ;
  END
END LUT4AB
END LIBRARY

