VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO N_term_single
  CLASS BLOCK ;
  FOREIGN N_term_single ;
  ORIGIN 0.000 0.000 ;
  SIZE 230.000 BY 50.000 ;
  PIN Ci
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.510 0.000 173.790 0.800 ;
    END
  END Ci
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 174.890 0.000 175.170 0.800 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 188.690 0.000 188.970 0.800 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 190.070 0.000 190.350 0.800 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 191.450 0.000 191.730 0.800 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 192.830 0.000 193.110 0.800 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 194.210 0.000 194.490 0.800 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 195.590 0.000 195.870 0.800 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 196.970 0.000 197.250 0.800 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 198.350 0.000 198.630 0.800 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 0.800 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 201.110 0.000 201.390 0.800 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 176.270 0.000 176.550 0.800 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 177.650 0.000 177.930 0.800 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 179.030 0.000 179.310 0.800 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 0.800 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 181.790 0.000 182.070 0.800 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 183.170 0.000 183.450 0.800 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 184.550 0.000 184.830 0.800 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 185.930 0.000 186.210 0.800 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 187.310 0.000 187.590 0.800 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 7.910 49.200 8.190 50.000 ;
    END
  END FrameStrobe_O[0]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 44.710 49.200 44.990 50.000 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 48.390 49.200 48.670 50.000 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 52.070 49.200 52.350 50.000 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 55.750 49.200 56.030 50.000 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 59.430 49.200 59.710 50.000 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 63.110 49.200 63.390 50.000 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 66.790 49.200 67.070 50.000 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 70.470 49.200 70.750 50.000 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 74.150 49.200 74.430 50.000 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 77.830 49.200 78.110 50.000 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 11.590 49.200 11.870 50.000 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 15.270 49.200 15.550 50.000 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 18.950 49.200 19.230 50.000 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 22.630 49.200 22.910 50.000 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 26.310 49.200 26.590 50.000 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 29.990 49.200 30.270 50.000 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 33.670 49.200 33.950 50.000 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 37.350 49.200 37.630 50.000 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 41.030 49.200 41.310 50.000 ;
    END
  END FrameStrobe_O[9]
  PIN N1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 28.610 0.000 28.890 0.800 ;
    END
  END N1END[0]
  PIN N1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 29.990 0.000 30.270 0.800 ;
    END
  END N1END[1]
  PIN N1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 31.370 0.000 31.650 0.800 ;
    END
  END N1END[2]
  PIN N1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 32.750 0.000 33.030 0.800 ;
    END
  END N1END[3]
  PIN N2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 0.800 ;
    END
  END N2END[0]
  PIN N2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 46.550 0.000 46.830 0.800 ;
    END
  END N2END[1]
  PIN N2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 47.930 0.000 48.210 0.800 ;
    END
  END N2END[2]
  PIN N2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 49.310 0.000 49.590 0.800 ;
    END
  END N2END[3]
  PIN N2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 50.690 0.000 50.970 0.800 ;
    END
  END N2END[4]
  PIN N2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 52.070 0.000 52.350 0.800 ;
    END
  END N2END[5]
  PIN N2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 53.450 0.000 53.730 0.800 ;
    END
  END N2END[6]
  PIN N2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 0.800 ;
    END
  END N2END[7]
  PIN N2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 34.130 0.000 34.410 0.800 ;
    END
  END N2MID[0]
  PIN N2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 0.800 ;
    END
  END N2MID[1]
  PIN N2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 36.890 0.000 37.170 0.800 ;
    END
  END N2MID[2]
  PIN N2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 38.270 0.000 38.550 0.800 ;
    END
  END N2MID[3]
  PIN N2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 39.650 0.000 39.930 0.800 ;
    END
  END N2MID[4]
  PIN N2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 41.030 0.000 41.310 0.800 ;
    END
  END N2MID[5]
  PIN N2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 42.410 0.000 42.690 0.800 ;
    END
  END N2MID[6]
  PIN N2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 43.790 0.000 44.070 0.800 ;
    END
  END N2MID[7]
  PIN N4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 56.210 0.000 56.490 0.800 ;
    END
  END N4END[0]
  PIN N4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 70.010 0.000 70.290 0.800 ;
    END
  END N4END[10]
  PIN N4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 71.390 0.000 71.670 0.800 ;
    END
  END N4END[11]
  PIN N4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 0.000 73.050 0.800 ;
    END
  END N4END[12]
  PIN N4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 0.800 ;
    END
  END N4END[13]
  PIN N4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.530 0.000 75.810 0.800 ;
    END
  END N4END[14]
  PIN N4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.910 0.000 77.190 0.800 ;
    END
  END N4END[15]
  PIN N4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 57.590 0.000 57.870 0.800 ;
    END
  END N4END[1]
  PIN N4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 58.970 0.000 59.250 0.800 ;
    END
  END N4END[2]
  PIN N4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 60.350 0.000 60.630 0.800 ;
    END
  END N4END[3]
  PIN N4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 61.730 0.000 62.010 0.800 ;
    END
  END N4END[4]
  PIN N4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 63.110 0.000 63.390 0.800 ;
    END
  END N4END[5]
  PIN N4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 0.800 ;
    END
  END N4END[6]
  PIN N4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 65.870 0.000 66.150 0.800 ;
    END
  END N4END[7]
  PIN N4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 67.250 0.000 67.530 0.800 ;
    END
  END N4END[8]
  PIN N4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 68.630 0.000 68.910 0.800 ;
    END
  END N4END[9]
  PIN NN4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 78.290 0.000 78.570 0.800 ;
    END
  END NN4END[0]
  PIN NN4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 92.090 0.000 92.370 0.800 ;
    END
  END NN4END[10]
  PIN NN4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 0.800 ;
    END
  END NN4END[11]
  PIN NN4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 94.850 0.000 95.130 0.800 ;
    END
  END NN4END[12]
  PIN NN4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 96.230 0.000 96.510 0.800 ;
    END
  END NN4END[13]
  PIN NN4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 97.610 0.000 97.890 0.800 ;
    END
  END NN4END[14]
  PIN NN4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 98.990 0.000 99.270 0.800 ;
    END
  END NN4END[15]
  PIN NN4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 79.670 0.000 79.950 0.800 ;
    END
  END NN4END[1]
  PIN NN4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 81.050 0.000 81.330 0.800 ;
    END
  END NN4END[2]
  PIN NN4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 82.430 0.000 82.710 0.800 ;
    END
  END NN4END[3]
  PIN NN4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 0.800 ;
    END
  END NN4END[4]
  PIN NN4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 85.190 0.000 85.470 0.800 ;
    END
  END NN4END[5]
  PIN NN4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 86.570 0.000 86.850 0.800 ;
    END
  END NN4END[6]
  PIN NN4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 87.950 0.000 88.230 0.800 ;
    END
  END NN4END[7]
  PIN NN4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 89.330 0.000 89.610 0.800 ;
    END
  END NN4END[8]
  PIN NN4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 90.710 0.000 90.990 0.800 ;
    END
  END NN4END[9]
  PIN S1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 100.370 0.000 100.650 0.800 ;
    END
  END S1BEG[0]
  PIN S1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 101.750 0.000 102.030 0.800 ;
    END
  END S1BEG[1]
  PIN S1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 0.800 ;
    END
  END S1BEG[2]
  PIN S1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 104.510 0.000 104.790 0.800 ;
    END
  END S1BEG[3]
  PIN S2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 116.930 0.000 117.210 0.800 ;
    END
  END S2BEG[0]
  PIN S2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 118.310 0.000 118.590 0.800 ;
    END
  END S2BEG[1]
  PIN S2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 0.800 ;
    END
  END S2BEG[2]
  PIN S2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 121.070 0.000 121.350 0.800 ;
    END
  END S2BEG[3]
  PIN S2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 0.800 ;
    END
  END S2BEG[4]
  PIN S2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 123.830 0.000 124.110 0.800 ;
    END
  END S2BEG[5]
  PIN S2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 125.210 0.000 125.490 0.800 ;
    END
  END S2BEG[6]
  PIN S2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 126.590 0.000 126.870 0.800 ;
    END
  END S2BEG[7]
  PIN S2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 105.890 0.000 106.170 0.800 ;
    END
  END S2BEGb[0]
  PIN S2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 107.270 0.000 107.550 0.800 ;
    END
  END S2BEGb[1]
  PIN S2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 108.650 0.000 108.930 0.800 ;
    END
  END S2BEGb[2]
  PIN S2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 110.030 0.000 110.310 0.800 ;
    END
  END S2BEGb[3]
  PIN S2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 111.410 0.000 111.690 0.800 ;
    END
  END S2BEGb[4]
  PIN S2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 0.800 ;
    END
  END S2BEGb[5]
  PIN S2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 114.170 0.000 114.450 0.800 ;
    END
  END S2BEGb[6]
  PIN S2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 115.550 0.000 115.830 0.800 ;
    END
  END S2BEGb[7]
  PIN S4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 127.970 0.000 128.250 0.800 ;
    END
  END S4BEG[0]
  PIN S4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 0.800 ;
    END
  END S4BEG[10]
  PIN S4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 143.150 0.000 143.430 0.800 ;
    END
  END S4BEG[11]
  PIN S4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 144.530 0.000 144.810 0.800 ;
    END
  END S4BEG[12]
  PIN S4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 145.910 0.000 146.190 0.800 ;
    END
  END S4BEG[13]
  PIN S4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 147.290 0.000 147.570 0.800 ;
    END
  END S4BEG[14]
  PIN S4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 148.670 0.000 148.950 0.800 ;
    END
  END S4BEG[15]
  PIN S4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 129.350 0.000 129.630 0.800 ;
    END
  END S4BEG[1]
  PIN S4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 130.730 0.000 131.010 0.800 ;
    END
  END S4BEG[2]
  PIN S4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 0.800 ;
    END
  END S4BEG[3]
  PIN S4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 133.490 0.000 133.770 0.800 ;
    END
  END S4BEG[4]
  PIN S4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 134.870 0.000 135.150 0.800 ;
    END
  END S4BEG[5]
  PIN S4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 136.250 0.000 136.530 0.800 ;
    END
  END S4BEG[6]
  PIN S4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 137.630 0.000 137.910 0.800 ;
    END
  END S4BEG[7]
  PIN S4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 139.010 0.000 139.290 0.800 ;
    END
  END S4BEG[8]
  PIN S4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 140.390 0.000 140.670 0.800 ;
    END
  END S4BEG[9]
  PIN SS4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 150.050 0.000 150.330 0.800 ;
    END
  END SS4BEG[0]
  PIN SS4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 163.850 0.000 164.130 0.800 ;
    END
  END SS4BEG[10]
  PIN SS4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 165.230 0.000 165.510 0.800 ;
    END
  END SS4BEG[11]
  PIN SS4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 166.610 0.000 166.890 0.800 ;
    END
  END SS4BEG[12]
  PIN SS4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 167.990 0.000 168.270 0.800 ;
    END
  END SS4BEG[13]
  PIN SS4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 169.370 0.000 169.650 0.800 ;
    END
  END SS4BEG[14]
  PIN SS4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 0.800 ;
    END
  END SS4BEG[15]
  PIN SS4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 151.430 0.000 151.710 0.800 ;
    END
  END SS4BEG[1]
  PIN SS4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 152.810 0.000 153.090 0.800 ;
    END
  END SS4BEG[2]
  PIN SS4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 154.190 0.000 154.470 0.800 ;
    END
  END SS4BEG[3]
  PIN SS4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 155.570 0.000 155.850 0.800 ;
    END
  END SS4BEG[4]
  PIN SS4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 156.950 0.000 157.230 0.800 ;
    END
  END SS4BEG[5]
  PIN SS4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 158.330 0.000 158.610 0.800 ;
    END
  END SS4BEG[6]
  PIN SS4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 159.710 0.000 159.990 0.800 ;
    END
  END SS4BEG[7]
  PIN SS4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 0.800 ;
    END
  END SS4BEG[8]
  PIN SS4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 162.470 0.000 162.750 0.800 ;
    END
  END SS4BEG[9]
  PIN UIO_TOP_UIN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 81.510 49.200 81.790 50.000 ;
    END
  END UIO_TOP_UIN0
  PIN UIO_TOP_UIN1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 85.190 49.200 85.470 50.000 ;
    END
  END UIO_TOP_UIN1
  PIN UIO_TOP_UIN10
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 88.870 49.200 89.150 50.000 ;
    END
  END UIO_TOP_UIN10
  PIN UIO_TOP_UIN11
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 92.550 49.200 92.830 50.000 ;
    END
  END UIO_TOP_UIN11
  PIN UIO_TOP_UIN12
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 96.230 49.200 96.510 50.000 ;
    END
  END UIO_TOP_UIN12
  PIN UIO_TOP_UIN13
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 99.910 49.200 100.190 50.000 ;
    END
  END UIO_TOP_UIN13
  PIN UIO_TOP_UIN14
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 103.590 49.200 103.870 50.000 ;
    END
  END UIO_TOP_UIN14
  PIN UIO_TOP_UIN15
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 107.270 49.200 107.550 50.000 ;
    END
  END UIO_TOP_UIN15
  PIN UIO_TOP_UIN16
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 110.950 49.200 111.230 50.000 ;
    END
  END UIO_TOP_UIN16
  PIN UIO_TOP_UIN17
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 114.630 49.200 114.910 50.000 ;
    END
  END UIO_TOP_UIN17
  PIN UIO_TOP_UIN18
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 118.310 49.200 118.590 50.000 ;
    END
  END UIO_TOP_UIN18
  PIN UIO_TOP_UIN19
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 121.990 49.200 122.270 50.000 ;
    END
  END UIO_TOP_UIN19
  PIN UIO_TOP_UIN2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 125.670 49.200 125.950 50.000 ;
    END
  END UIO_TOP_UIN2
  PIN UIO_TOP_UIN3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 129.350 49.200 129.630 50.000 ;
    END
  END UIO_TOP_UIN3
  PIN UIO_TOP_UIN4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 133.030 49.200 133.310 50.000 ;
    END
  END UIO_TOP_UIN4
  PIN UIO_TOP_UIN5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 136.710 49.200 136.990 50.000 ;
    END
  END UIO_TOP_UIN5
  PIN UIO_TOP_UIN6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 140.390 49.200 140.670 50.000 ;
    END
  END UIO_TOP_UIN6
  PIN UIO_TOP_UIN7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 144.070 49.200 144.350 50.000 ;
    END
  END UIO_TOP_UIN7
  PIN UIO_TOP_UIN8
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 147.750 49.200 148.030 50.000 ;
    END
  END UIO_TOP_UIN8
  PIN UIO_TOP_UIN9
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 151.430 49.200 151.710 50.000 ;
    END
  END UIO_TOP_UIN9
  PIN UIO_TOP_UOUT0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 155.110 49.200 155.390 50.000 ;
    END
  END UIO_TOP_UOUT0
  PIN UIO_TOP_UOUT1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 158.790 49.200 159.070 50.000 ;
    END
  END UIO_TOP_UOUT1
  PIN UIO_TOP_UOUT10
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 162.470 49.200 162.750 50.000 ;
    END
  END UIO_TOP_UOUT10
  PIN UIO_TOP_UOUT11
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 166.150 49.200 166.430 50.000 ;
    END
  END UIO_TOP_UOUT11
  PIN UIO_TOP_UOUT12
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 169.830 49.200 170.110 50.000 ;
    END
  END UIO_TOP_UOUT12
  PIN UIO_TOP_UOUT13
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 173.510 49.200 173.790 50.000 ;
    END
  END UIO_TOP_UOUT13
  PIN UIO_TOP_UOUT14
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 177.190 49.200 177.470 50.000 ;
    END
  END UIO_TOP_UOUT14
  PIN UIO_TOP_UOUT15
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 180.870 49.200 181.150 50.000 ;
    END
  END UIO_TOP_UOUT15
  PIN UIO_TOP_UOUT16
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 184.550 49.200 184.830 50.000 ;
    END
  END UIO_TOP_UOUT16
  PIN UIO_TOP_UOUT17
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 188.230 49.200 188.510 50.000 ;
    END
  END UIO_TOP_UOUT17
  PIN UIO_TOP_UOUT18
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 191.910 49.200 192.190 50.000 ;
    END
  END UIO_TOP_UOUT18
  PIN UIO_TOP_UOUT19
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 195.590 49.200 195.870 50.000 ;
    END
  END UIO_TOP_UOUT19
  PIN UIO_TOP_UOUT2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 199.270 49.200 199.550 50.000 ;
    END
  END UIO_TOP_UOUT2
  PIN UIO_TOP_UOUT3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 202.950 49.200 203.230 50.000 ;
    END
  END UIO_TOP_UOUT3
  PIN UIO_TOP_UOUT4
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 206.630 49.200 206.910 50.000 ;
    END
  END UIO_TOP_UOUT4
  PIN UIO_TOP_UOUT5
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 210.310 49.200 210.590 50.000 ;
    END
  END UIO_TOP_UOUT5
  PIN UIO_TOP_UOUT6
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 213.990 49.200 214.270 50.000 ;
    END
  END UIO_TOP_UOUT6
  PIN UIO_TOP_UOUT7
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 217.670 49.200 217.950 50.000 ;
    END
  END UIO_TOP_UOUT7
  PIN UIO_TOP_UOUT8
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 221.350 49.200 221.630 50.000 ;
    END
  END UIO_TOP_UOUT8
  PIN UIO_TOP_UOUT9
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 225.030 49.200 225.310 50.000 ;
    END
  END UIO_TOP_UOUT9
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 172.130 0.000 172.410 0.800 ;
    END
  END UserCLK
  PIN UserCLKo
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 4.230 49.200 4.510 50.000 ;
    END
  END UserCLKo
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 32.085 10.640 33.685 38.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 86.820 10.640 88.420 38.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 141.555 10.640 143.155 38.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 196.290 10.640 197.890 38.320 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 59.450 10.640 61.050 38.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 114.185 10.640 115.785 38.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 168.920 10.640 170.520 38.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 223.655 10.640 225.255 38.320 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 224.480 38.165 ;
      LAYER met1 ;
        RECT 4.210 5.480 225.790 41.100 ;
      LAYER met2 ;
        RECT 4.790 48.920 7.630 49.370 ;
        RECT 8.470 48.920 11.310 49.370 ;
        RECT 12.150 48.920 14.990 49.370 ;
        RECT 15.830 48.920 18.670 49.370 ;
        RECT 19.510 48.920 22.350 49.370 ;
        RECT 23.190 48.920 26.030 49.370 ;
        RECT 26.870 48.920 29.710 49.370 ;
        RECT 30.550 48.920 33.390 49.370 ;
        RECT 34.230 48.920 37.070 49.370 ;
        RECT 37.910 48.920 40.750 49.370 ;
        RECT 41.590 48.920 44.430 49.370 ;
        RECT 45.270 48.920 48.110 49.370 ;
        RECT 48.950 48.920 51.790 49.370 ;
        RECT 52.630 48.920 55.470 49.370 ;
        RECT 56.310 48.920 59.150 49.370 ;
        RECT 59.990 48.920 62.830 49.370 ;
        RECT 63.670 48.920 66.510 49.370 ;
        RECT 67.350 48.920 70.190 49.370 ;
        RECT 71.030 48.920 73.870 49.370 ;
        RECT 74.710 48.920 77.550 49.370 ;
        RECT 78.390 48.920 81.230 49.370 ;
        RECT 82.070 48.920 84.910 49.370 ;
        RECT 85.750 48.920 88.590 49.370 ;
        RECT 89.430 48.920 92.270 49.370 ;
        RECT 93.110 48.920 95.950 49.370 ;
        RECT 96.790 48.920 99.630 49.370 ;
        RECT 100.470 48.920 103.310 49.370 ;
        RECT 104.150 48.920 106.990 49.370 ;
        RECT 107.830 48.920 110.670 49.370 ;
        RECT 111.510 48.920 114.350 49.370 ;
        RECT 115.190 48.920 118.030 49.370 ;
        RECT 118.870 48.920 121.710 49.370 ;
        RECT 122.550 48.920 125.390 49.370 ;
        RECT 126.230 48.920 129.070 49.370 ;
        RECT 129.910 48.920 132.750 49.370 ;
        RECT 133.590 48.920 136.430 49.370 ;
        RECT 137.270 48.920 140.110 49.370 ;
        RECT 140.950 48.920 143.790 49.370 ;
        RECT 144.630 48.920 147.470 49.370 ;
        RECT 148.310 48.920 151.150 49.370 ;
        RECT 151.990 48.920 154.830 49.370 ;
        RECT 155.670 48.920 158.510 49.370 ;
        RECT 159.350 48.920 162.190 49.370 ;
        RECT 163.030 48.920 165.870 49.370 ;
        RECT 166.710 48.920 169.550 49.370 ;
        RECT 170.390 48.920 173.230 49.370 ;
        RECT 174.070 48.920 176.910 49.370 ;
        RECT 177.750 48.920 180.590 49.370 ;
        RECT 181.430 48.920 184.270 49.370 ;
        RECT 185.110 48.920 187.950 49.370 ;
        RECT 188.790 48.920 191.630 49.370 ;
        RECT 192.470 48.920 195.310 49.370 ;
        RECT 196.150 48.920 198.990 49.370 ;
        RECT 199.830 48.920 202.670 49.370 ;
        RECT 203.510 48.920 206.350 49.370 ;
        RECT 207.190 48.920 210.030 49.370 ;
        RECT 210.870 48.920 213.710 49.370 ;
        RECT 214.550 48.920 217.390 49.370 ;
        RECT 218.230 48.920 221.070 49.370 ;
        RECT 221.910 48.920 224.750 49.370 ;
        RECT 225.590 48.920 225.760 49.370 ;
        RECT 4.240 1.080 225.760 48.920 ;
        RECT 4.240 0.155 28.330 1.080 ;
        RECT 29.170 0.155 29.710 1.080 ;
        RECT 30.550 0.155 31.090 1.080 ;
        RECT 31.930 0.155 32.470 1.080 ;
        RECT 33.310 0.155 33.850 1.080 ;
        RECT 34.690 0.155 35.230 1.080 ;
        RECT 36.070 0.155 36.610 1.080 ;
        RECT 37.450 0.155 37.990 1.080 ;
        RECT 38.830 0.155 39.370 1.080 ;
        RECT 40.210 0.155 40.750 1.080 ;
        RECT 41.590 0.155 42.130 1.080 ;
        RECT 42.970 0.155 43.510 1.080 ;
        RECT 44.350 0.155 44.890 1.080 ;
        RECT 45.730 0.155 46.270 1.080 ;
        RECT 47.110 0.155 47.650 1.080 ;
        RECT 48.490 0.155 49.030 1.080 ;
        RECT 49.870 0.155 50.410 1.080 ;
        RECT 51.250 0.155 51.790 1.080 ;
        RECT 52.630 0.155 53.170 1.080 ;
        RECT 54.010 0.155 54.550 1.080 ;
        RECT 55.390 0.155 55.930 1.080 ;
        RECT 56.770 0.155 57.310 1.080 ;
        RECT 58.150 0.155 58.690 1.080 ;
        RECT 59.530 0.155 60.070 1.080 ;
        RECT 60.910 0.155 61.450 1.080 ;
        RECT 62.290 0.155 62.830 1.080 ;
        RECT 63.670 0.155 64.210 1.080 ;
        RECT 65.050 0.155 65.590 1.080 ;
        RECT 66.430 0.155 66.970 1.080 ;
        RECT 67.810 0.155 68.350 1.080 ;
        RECT 69.190 0.155 69.730 1.080 ;
        RECT 70.570 0.155 71.110 1.080 ;
        RECT 71.950 0.155 72.490 1.080 ;
        RECT 73.330 0.155 73.870 1.080 ;
        RECT 74.710 0.155 75.250 1.080 ;
        RECT 76.090 0.155 76.630 1.080 ;
        RECT 77.470 0.155 78.010 1.080 ;
        RECT 78.850 0.155 79.390 1.080 ;
        RECT 80.230 0.155 80.770 1.080 ;
        RECT 81.610 0.155 82.150 1.080 ;
        RECT 82.990 0.155 83.530 1.080 ;
        RECT 84.370 0.155 84.910 1.080 ;
        RECT 85.750 0.155 86.290 1.080 ;
        RECT 87.130 0.155 87.670 1.080 ;
        RECT 88.510 0.155 89.050 1.080 ;
        RECT 89.890 0.155 90.430 1.080 ;
        RECT 91.270 0.155 91.810 1.080 ;
        RECT 92.650 0.155 93.190 1.080 ;
        RECT 94.030 0.155 94.570 1.080 ;
        RECT 95.410 0.155 95.950 1.080 ;
        RECT 96.790 0.155 97.330 1.080 ;
        RECT 98.170 0.155 98.710 1.080 ;
        RECT 99.550 0.155 100.090 1.080 ;
        RECT 100.930 0.155 101.470 1.080 ;
        RECT 102.310 0.155 102.850 1.080 ;
        RECT 103.690 0.155 104.230 1.080 ;
        RECT 105.070 0.155 105.610 1.080 ;
        RECT 106.450 0.155 106.990 1.080 ;
        RECT 107.830 0.155 108.370 1.080 ;
        RECT 109.210 0.155 109.750 1.080 ;
        RECT 110.590 0.155 111.130 1.080 ;
        RECT 111.970 0.155 112.510 1.080 ;
        RECT 113.350 0.155 113.890 1.080 ;
        RECT 114.730 0.155 115.270 1.080 ;
        RECT 116.110 0.155 116.650 1.080 ;
        RECT 117.490 0.155 118.030 1.080 ;
        RECT 118.870 0.155 119.410 1.080 ;
        RECT 120.250 0.155 120.790 1.080 ;
        RECT 121.630 0.155 122.170 1.080 ;
        RECT 123.010 0.155 123.550 1.080 ;
        RECT 124.390 0.155 124.930 1.080 ;
        RECT 125.770 0.155 126.310 1.080 ;
        RECT 127.150 0.155 127.690 1.080 ;
        RECT 128.530 0.155 129.070 1.080 ;
        RECT 129.910 0.155 130.450 1.080 ;
        RECT 131.290 0.155 131.830 1.080 ;
        RECT 132.670 0.155 133.210 1.080 ;
        RECT 134.050 0.155 134.590 1.080 ;
        RECT 135.430 0.155 135.970 1.080 ;
        RECT 136.810 0.155 137.350 1.080 ;
        RECT 138.190 0.155 138.730 1.080 ;
        RECT 139.570 0.155 140.110 1.080 ;
        RECT 140.950 0.155 141.490 1.080 ;
        RECT 142.330 0.155 142.870 1.080 ;
        RECT 143.710 0.155 144.250 1.080 ;
        RECT 145.090 0.155 145.630 1.080 ;
        RECT 146.470 0.155 147.010 1.080 ;
        RECT 147.850 0.155 148.390 1.080 ;
        RECT 149.230 0.155 149.770 1.080 ;
        RECT 150.610 0.155 151.150 1.080 ;
        RECT 151.990 0.155 152.530 1.080 ;
        RECT 153.370 0.155 153.910 1.080 ;
        RECT 154.750 0.155 155.290 1.080 ;
        RECT 156.130 0.155 156.670 1.080 ;
        RECT 157.510 0.155 158.050 1.080 ;
        RECT 158.890 0.155 159.430 1.080 ;
        RECT 160.270 0.155 160.810 1.080 ;
        RECT 161.650 0.155 162.190 1.080 ;
        RECT 163.030 0.155 163.570 1.080 ;
        RECT 164.410 0.155 164.950 1.080 ;
        RECT 165.790 0.155 166.330 1.080 ;
        RECT 167.170 0.155 167.710 1.080 ;
        RECT 168.550 0.155 169.090 1.080 ;
        RECT 169.930 0.155 170.470 1.080 ;
        RECT 171.310 0.155 171.850 1.080 ;
        RECT 172.690 0.155 173.230 1.080 ;
        RECT 174.070 0.155 174.610 1.080 ;
        RECT 175.450 0.155 175.990 1.080 ;
        RECT 176.830 0.155 177.370 1.080 ;
        RECT 178.210 0.155 178.750 1.080 ;
        RECT 179.590 0.155 180.130 1.080 ;
        RECT 180.970 0.155 181.510 1.080 ;
        RECT 182.350 0.155 182.890 1.080 ;
        RECT 183.730 0.155 184.270 1.080 ;
        RECT 185.110 0.155 185.650 1.080 ;
        RECT 186.490 0.155 187.030 1.080 ;
        RECT 187.870 0.155 188.410 1.080 ;
        RECT 189.250 0.155 189.790 1.080 ;
        RECT 190.630 0.155 191.170 1.080 ;
        RECT 192.010 0.155 192.550 1.080 ;
        RECT 193.390 0.155 193.930 1.080 ;
        RECT 194.770 0.155 195.310 1.080 ;
        RECT 196.150 0.155 196.690 1.080 ;
        RECT 197.530 0.155 198.070 1.080 ;
        RECT 198.910 0.155 199.450 1.080 ;
        RECT 200.290 0.155 200.830 1.080 ;
        RECT 201.670 0.155 225.760 1.080 ;
      LAYER met3 ;
        RECT 8.805 0.175 225.245 39.945 ;
      LAYER met4 ;
        RECT 94.135 10.240 113.785 21.585 ;
        RECT 116.185 10.240 141.155 21.585 ;
        RECT 143.555 10.240 159.785 21.585 ;
        RECT 94.135 0.175 159.785 10.240 ;
  END
END N_term_single
END LIBRARY

