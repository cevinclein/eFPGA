VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO RAM_IO
  CLASS BLOCK ;
  FOREIGN RAM_IO ;
  ORIGIN 0.000 0.000 ;
  SIZE 130.000 BY 223.115 ;
  PIN Config_accessC_bit0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 129.200 46.280 130.000 46.880 ;
    END
  END Config_accessC_bit0
  PIN Config_accessC_bit1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 129.200 49.000 130.000 49.600 ;
    END
  END Config_accessC_bit1
  PIN Config_accessC_bit2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 129.200 51.720 130.000 52.320 ;
    END
  END Config_accessC_bit2
  PIN Config_accessC_bit3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 129.200 54.440 130.000 55.040 ;
    END
  END Config_accessC_bit3
  PIN E1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 0.800 90.400 ;
    END
  END E1END[0]
  PIN E1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 0.800 91.760 ;
    END
  END E1END[1]
  PIN E1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 0.800 93.120 ;
    END
  END E1END[2]
  PIN E1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 0.800 94.480 ;
    END
  END E1END[3]
  PIN E2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.120 0.800 106.720 ;
    END
  END E2END[0]
  PIN E2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 0.800 108.080 ;
    END
  END E2END[1]
  PIN E2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 0.800 109.440 ;
    END
  END E2END[2]
  PIN E2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 0.800 110.800 ;
    END
  END E2END[3]
  PIN E2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.560 0.800 112.160 ;
    END
  END E2END[4]
  PIN E2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 0.800 113.520 ;
    END
  END E2END[5]
  PIN E2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.280 0.800 114.880 ;
    END
  END E2END[6]
  PIN E2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 0.800 116.240 ;
    END
  END E2END[7]
  PIN E2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 0.800 95.840 ;
    END
  END E2MID[0]
  PIN E2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 0.800 97.200 ;
    END
  END E2MID[1]
  PIN E2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 0.800 98.560 ;
    END
  END E2MID[2]
  PIN E2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.320 0.800 99.920 ;
    END
  END E2MID[3]
  PIN E2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 0.800 101.280 ;
    END
  END E2MID[4]
  PIN E2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 0.800 102.640 ;
    END
  END E2MID[5]
  PIN E2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 0.800 104.000 ;
    END
  END E2MID[6]
  PIN E2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.760 0.800 105.360 ;
    END
  END E2MID[7]
  PIN E6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.760 0.800 139.360 ;
    END
  END E6END[0]
  PIN E6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.360 0.800 152.960 ;
    END
  END E6END[10]
  PIN E6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.720 0.800 154.320 ;
    END
  END E6END[11]
  PIN E6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.120 0.800 140.720 ;
    END
  END E6END[1]
  PIN E6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.480 0.800 142.080 ;
    END
  END E6END[2]
  PIN E6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 0.800 143.440 ;
    END
  END E6END[3]
  PIN E6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.200 0.800 144.800 ;
    END
  END E6END[4]
  PIN E6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 0.800 146.160 ;
    END
  END E6END[5]
  PIN E6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.920 0.800 147.520 ;
    END
  END E6END[6]
  PIN E6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.280 0.800 148.880 ;
    END
  END E6END[7]
  PIN E6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 0.800 150.240 ;
    END
  END E6END[8]
  PIN E6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.000 0.800 151.600 ;
    END
  END E6END[9]
  PIN EE4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 0.800 117.600 ;
    END
  END EE4END[0]
  PIN EE4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 0.800 131.200 ;
    END
  END EE4END[10]
  PIN EE4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.960 0.800 132.560 ;
    END
  END EE4END[11]
  PIN EE4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.320 0.800 133.920 ;
    END
  END EE4END[12]
  PIN EE4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.680 0.800 135.280 ;
    END
  END EE4END[13]
  PIN EE4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 0.800 136.640 ;
    END
  END EE4END[14]
  PIN EE4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 0.800 138.000 ;
    END
  END EE4END[15]
  PIN EE4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.360 0.800 118.960 ;
    END
  END EE4END[1]
  PIN EE4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 0.800 120.320 ;
    END
  END EE4END[2]
  PIN EE4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 0.800 121.680 ;
    END
  END EE4END[3]
  PIN EE4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 0.800 123.040 ;
    END
  END EE4END[4]
  PIN EE4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.800 0.800 124.400 ;
    END
  END EE4END[5]
  PIN EE4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.160 0.800 125.760 ;
    END
  END EE4END[6]
  PIN EE4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 0.800 127.120 ;
    END
  END EE4END[7]
  PIN EE4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 0.800 128.480 ;
    END
  END EE4END[8]
  PIN EE4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 0.800 129.840 ;
    END
  END EE4END[9]
  PIN FAB2RAM_A0_O0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 129.200 78.920 130.000 79.520 ;
    END
  END FAB2RAM_A0_O0
  PIN FAB2RAM_A0_O1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 129.200 81.640 130.000 82.240 ;
    END
  END FAB2RAM_A0_O1
  PIN FAB2RAM_A0_O2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 129.200 84.360 130.000 84.960 ;
    END
  END FAB2RAM_A0_O2
  PIN FAB2RAM_A0_O3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 129.200 87.080 130.000 87.680 ;
    END
  END FAB2RAM_A0_O3
  PIN FAB2RAM_A1_O0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 129.200 68.040 130.000 68.640 ;
    END
  END FAB2RAM_A1_O0
  PIN FAB2RAM_A1_O1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 129.200 70.760 130.000 71.360 ;
    END
  END FAB2RAM_A1_O1
  PIN FAB2RAM_A1_O2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 129.200 73.480 130.000 74.080 ;
    END
  END FAB2RAM_A1_O2
  PIN FAB2RAM_A1_O3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 129.200 76.200 130.000 76.800 ;
    END
  END FAB2RAM_A1_O3
  PIN FAB2RAM_C_O0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 129.200 57.160 130.000 57.760 ;
    END
  END FAB2RAM_C_O0
  PIN FAB2RAM_C_O1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 129.200 59.880 130.000 60.480 ;
    END
  END FAB2RAM_C_O1
  PIN FAB2RAM_C_O2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 129.200 62.600 130.000 63.200 ;
    END
  END FAB2RAM_C_O2
  PIN FAB2RAM_C_O3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 129.200 65.320 130.000 65.920 ;
    END
  END FAB2RAM_C_O3
  PIN FAB2RAM_D0_O0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 129.200 122.440 130.000 123.040 ;
    END
  END FAB2RAM_D0_O0
  PIN FAB2RAM_D0_O1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 129.200 125.160 130.000 125.760 ;
    END
  END FAB2RAM_D0_O1
  PIN FAB2RAM_D0_O2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 129.200 127.880 130.000 128.480 ;
    END
  END FAB2RAM_D0_O2
  PIN FAB2RAM_D0_O3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 129.200 130.600 130.000 131.200 ;
    END
  END FAB2RAM_D0_O3
  PIN FAB2RAM_D1_O0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 129.200 111.560 130.000 112.160 ;
    END
  END FAB2RAM_D1_O0
  PIN FAB2RAM_D1_O1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 129.200 114.280 130.000 114.880 ;
    END
  END FAB2RAM_D1_O1
  PIN FAB2RAM_D1_O2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 129.200 117.000 130.000 117.600 ;
    END
  END FAB2RAM_D1_O2
  PIN FAB2RAM_D1_O3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 129.200 119.720 130.000 120.320 ;
    END
  END FAB2RAM_D1_O3
  PIN FAB2RAM_D2_O0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 129.200 100.680 130.000 101.280 ;
    END
  END FAB2RAM_D2_O0
  PIN FAB2RAM_D2_O1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 129.200 103.400 130.000 104.000 ;
    END
  END FAB2RAM_D2_O1
  PIN FAB2RAM_D2_O2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 129.200 106.120 130.000 106.720 ;
    END
  END FAB2RAM_D2_O2
  PIN FAB2RAM_D2_O3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 129.200 108.840 130.000 109.440 ;
    END
  END FAB2RAM_D2_O3
  PIN FAB2RAM_D3_O0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 129.200 89.800 130.000 90.400 ;
    END
  END FAB2RAM_D3_O0
  PIN FAB2RAM_D3_O1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 129.200 92.520 130.000 93.120 ;
    END
  END FAB2RAM_D3_O1
  PIN FAB2RAM_D3_O2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 129.200 95.240 130.000 95.840 ;
    END
  END FAB2RAM_D3_O2
  PIN FAB2RAM_D3_O3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 129.200 97.960 130.000 98.560 ;
    END
  END FAB2RAM_D3_O3
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.080 0.800 155.680 ;
    END
  END FrameData[0]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.680 0.800 169.280 ;
    END
  END FrameData[10]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 0.800 170.640 ;
    END
  END FrameData[11]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 171.400 0.800 172.000 ;
    END
  END FrameData[12]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.760 0.800 173.360 ;
    END
  END FrameData[13]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.120 0.800 174.720 ;
    END
  END FrameData[14]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.480 0.800 176.080 ;
    END
  END FrameData[15]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 0.800 177.440 ;
    END
  END FrameData[16]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.200 0.800 178.800 ;
    END
  END FrameData[17]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.560 0.800 180.160 ;
    END
  END FrameData[18]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.920 0.800 181.520 ;
    END
  END FrameData[19]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 0.800 157.040 ;
    END
  END FrameData[1]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.280 0.800 182.880 ;
    END
  END FrameData[20]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 0.800 184.240 ;
    END
  END FrameData[21]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.000 0.800 185.600 ;
    END
  END FrameData[22]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 186.360 0.800 186.960 ;
    END
  END FrameData[23]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.720 0.800 188.320 ;
    END
  END FrameData[24]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.080 0.800 189.680 ;
    END
  END FrameData[25]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 0.800 191.040 ;
    END
  END FrameData[26]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.800 0.800 192.400 ;
    END
  END FrameData[27]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 0.800 193.760 ;
    END
  END FrameData[28]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 194.520 0.800 195.120 ;
    END
  END FrameData[29]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.800 0.800 158.400 ;
    END
  END FrameData[2]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.880 0.800 196.480 ;
    END
  END FrameData[30]
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 0.800 197.840 ;
    END
  END FrameData[31]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.160 0.800 159.760 ;
    END
  END FrameData[3]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.520 0.800 161.120 ;
    END
  END FrameData[4]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.880 0.800 162.480 ;
    END
  END FrameData[5]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 0.800 163.840 ;
    END
  END FrameData[6]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.600 0.800 165.200 ;
    END
  END FrameData[7]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.960 0.800 166.560 ;
    END
  END FrameData[8]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 167.320 0.800 167.920 ;
    END
  END FrameData[9]
  PIN FrameData_O[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 129.200 133.320 130.000 133.920 ;
    END
  END FrameData_O[0]
  PIN FrameData_O[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 129.200 160.520 130.000 161.120 ;
    END
  END FrameData_O[10]
  PIN FrameData_O[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 129.200 163.240 130.000 163.840 ;
    END
  END FrameData_O[11]
  PIN FrameData_O[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 129.200 165.960 130.000 166.560 ;
    END
  END FrameData_O[12]
  PIN FrameData_O[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 129.200 168.680 130.000 169.280 ;
    END
  END FrameData_O[13]
  PIN FrameData_O[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 129.200 171.400 130.000 172.000 ;
    END
  END FrameData_O[14]
  PIN FrameData_O[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 129.200 174.120 130.000 174.720 ;
    END
  END FrameData_O[15]
  PIN FrameData_O[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 129.200 176.840 130.000 177.440 ;
    END
  END FrameData_O[16]
  PIN FrameData_O[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 129.200 179.560 130.000 180.160 ;
    END
  END FrameData_O[17]
  PIN FrameData_O[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 129.200 182.280 130.000 182.880 ;
    END
  END FrameData_O[18]
  PIN FrameData_O[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 129.200 185.000 130.000 185.600 ;
    END
  END FrameData_O[19]
  PIN FrameData_O[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 129.200 136.040 130.000 136.640 ;
    END
  END FrameData_O[1]
  PIN FrameData_O[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 129.200 187.720 130.000 188.320 ;
    END
  END FrameData_O[20]
  PIN FrameData_O[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 129.200 190.440 130.000 191.040 ;
    END
  END FrameData_O[21]
  PIN FrameData_O[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 129.200 193.160 130.000 193.760 ;
    END
  END FrameData_O[22]
  PIN FrameData_O[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 129.200 195.880 130.000 196.480 ;
    END
  END FrameData_O[23]
  PIN FrameData_O[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 129.200 198.600 130.000 199.200 ;
    END
  END FrameData_O[24]
  PIN FrameData_O[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 129.200 201.320 130.000 201.920 ;
    END
  END FrameData_O[25]
  PIN FrameData_O[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 129.200 204.040 130.000 204.640 ;
    END
  END FrameData_O[26]
  PIN FrameData_O[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 129.200 206.760 130.000 207.360 ;
    END
  END FrameData_O[27]
  PIN FrameData_O[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 129.200 209.480 130.000 210.080 ;
    END
  END FrameData_O[28]
  PIN FrameData_O[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 129.200 212.200 130.000 212.800 ;
    END
  END FrameData_O[29]
  PIN FrameData_O[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 129.200 138.760 130.000 139.360 ;
    END
  END FrameData_O[2]
  PIN FrameData_O[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 129.200 214.920 130.000 215.520 ;
    END
  END FrameData_O[30]
  PIN FrameData_O[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 129.200 217.640 130.000 218.240 ;
    END
  END FrameData_O[31]
  PIN FrameData_O[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 129.200 141.480 130.000 142.080 ;
    END
  END FrameData_O[3]
  PIN FrameData_O[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 129.200 144.200 130.000 144.800 ;
    END
  END FrameData_O[4]
  PIN FrameData_O[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 129.200 146.920 130.000 147.520 ;
    END
  END FrameData_O[5]
  PIN FrameData_O[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 129.200 149.640 130.000 150.240 ;
    END
  END FrameData_O[6]
  PIN FrameData_O[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 129.200 152.360 130.000 152.960 ;
    END
  END FrameData_O[7]
  PIN FrameData_O[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 129.200 155.080 130.000 155.680 ;
    END
  END FrameData_O[8]
  PIN FrameData_O[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 129.200 157.800 130.000 158.400 ;
    END
  END FrameData_O[9]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 101.750 0.000 102.030 0.800 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 115.550 0.000 115.830 0.800 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 116.930 0.000 117.210 0.800 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 118.310 0.000 118.590 0.800 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 0.800 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 121.070 0.000 121.350 0.800 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 0.800 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 123.830 0.000 124.110 0.800 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 125.210 0.000 125.490 0.800 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 126.590 0.000 126.870 0.800 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 127.970 0.000 128.250 0.800 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 0.800 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 104.510 0.000 104.790 0.800 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 105.890 0.000 106.170 0.800 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 107.270 0.000 107.550 0.800 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 108.650 0.000 108.930 0.800 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 110.030 0.000 110.310 0.800 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 111.410 0.000 111.690 0.800 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 0.800 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 114.170 0.000 114.450 0.800 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 101.750 222.315 102.030 223.115 ;
    END
  END FrameStrobe_O[0]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 115.550 222.315 115.830 223.115 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 116.930 222.315 117.210 223.115 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 118.310 222.315 118.590 223.115 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 119.690 222.315 119.970 223.115 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 121.070 222.315 121.350 223.115 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 122.450 222.315 122.730 223.115 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 123.830 222.315 124.110 223.115 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 125.210 222.315 125.490 223.115 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 126.590 222.315 126.870 223.115 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 127.970 222.315 128.250 223.115 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 103.130 222.315 103.410 223.115 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 104.510 222.315 104.790 223.115 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 105.890 222.315 106.170 223.115 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 107.270 222.315 107.550 223.115 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 108.650 222.315 108.930 223.115 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 110.030 222.315 110.310 223.115 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 111.410 222.315 111.690 223.115 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 112.790 222.315 113.070 223.115 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 114.170 222.315 114.450 223.115 ;
    END
  END FrameStrobe_O[9]
  PIN N1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 1.010 222.315 1.290 223.115 ;
    END
  END N1BEG[0]
  PIN N1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 2.390 222.315 2.670 223.115 ;
    END
  END N1BEG[1]
  PIN N1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 3.770 222.315 4.050 223.115 ;
    END
  END N1BEG[2]
  PIN N1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 5.150 222.315 5.430 223.115 ;
    END
  END N1BEG[3]
  PIN N1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 1.010 0.000 1.290 0.800 ;
    END
  END N1END[0]
  PIN N1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 2.390 0.000 2.670 0.800 ;
    END
  END N1END[1]
  PIN N1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 3.770 0.000 4.050 0.800 ;
    END
  END N1END[2]
  PIN N1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 5.150 0.000 5.430 0.800 ;
    END
  END N1END[3]
  PIN N2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 6.530 222.315 6.810 223.115 ;
    END
  END N2BEG[0]
  PIN N2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 7.910 222.315 8.190 223.115 ;
    END
  END N2BEG[1]
  PIN N2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 9.290 222.315 9.570 223.115 ;
    END
  END N2BEG[2]
  PIN N2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 10.670 222.315 10.950 223.115 ;
    END
  END N2BEG[3]
  PIN N2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 12.050 222.315 12.330 223.115 ;
    END
  END N2BEG[4]
  PIN N2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 13.430 222.315 13.710 223.115 ;
    END
  END N2BEG[5]
  PIN N2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 14.810 222.315 15.090 223.115 ;
    END
  END N2BEG[6]
  PIN N2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 16.190 222.315 16.470 223.115 ;
    END
  END N2BEG[7]
  PIN N2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 17.570 222.315 17.850 223.115 ;
    END
  END N2BEGb[0]
  PIN N2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 18.950 222.315 19.230 223.115 ;
    END
  END N2BEGb[1]
  PIN N2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 20.330 222.315 20.610 223.115 ;
    END
  END N2BEGb[2]
  PIN N2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 21.710 222.315 21.990 223.115 ;
    END
  END N2BEGb[3]
  PIN N2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 23.090 222.315 23.370 223.115 ;
    END
  END N2BEGb[4]
  PIN N2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 24.470 222.315 24.750 223.115 ;
    END
  END N2BEGb[5]
  PIN N2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 25.850 222.315 26.130 223.115 ;
    END
  END N2BEGb[6]
  PIN N2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 27.230 222.315 27.510 223.115 ;
    END
  END N2BEGb[7]
  PIN N2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 17.570 0.000 17.850 0.800 ;
    END
  END N2END[0]
  PIN N2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 18.950 0.000 19.230 0.800 ;
    END
  END N2END[1]
  PIN N2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 20.330 0.000 20.610 0.800 ;
    END
  END N2END[2]
  PIN N2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 21.710 0.000 21.990 0.800 ;
    END
  END N2END[3]
  PIN N2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 23.090 0.000 23.370 0.800 ;
    END
  END N2END[4]
  PIN N2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 24.470 0.000 24.750 0.800 ;
    END
  END N2END[5]
  PIN N2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 0.800 ;
    END
  END N2END[6]
  PIN N2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 27.230 0.000 27.510 0.800 ;
    END
  END N2END[7]
  PIN N2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 0.800 ;
    END
  END N2MID[0]
  PIN N2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 7.910 0.000 8.190 0.800 ;
    END
  END N2MID[1]
  PIN N2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 9.290 0.000 9.570 0.800 ;
    END
  END N2MID[2]
  PIN N2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 10.670 0.000 10.950 0.800 ;
    END
  END N2MID[3]
  PIN N2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 12.050 0.000 12.330 0.800 ;
    END
  END N2MID[4]
  PIN N2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 13.430 0.000 13.710 0.800 ;
    END
  END N2MID[5]
  PIN N2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 14.810 0.000 15.090 0.800 ;
    END
  END N2MID[6]
  PIN N2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 0.800 ;
    END
  END N2MID[7]
  PIN N4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 28.610 222.315 28.890 223.115 ;
    END
  END N4BEG[0]
  PIN N4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 42.410 222.315 42.690 223.115 ;
    END
  END N4BEG[10]
  PIN N4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 43.790 222.315 44.070 223.115 ;
    END
  END N4BEG[11]
  PIN N4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 45.170 222.315 45.450 223.115 ;
    END
  END N4BEG[12]
  PIN N4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 46.550 222.315 46.830 223.115 ;
    END
  END N4BEG[13]
  PIN N4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 47.930 222.315 48.210 223.115 ;
    END
  END N4BEG[14]
  PIN N4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 49.310 222.315 49.590 223.115 ;
    END
  END N4BEG[15]
  PIN N4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 29.990 222.315 30.270 223.115 ;
    END
  END N4BEG[1]
  PIN N4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 31.370 222.315 31.650 223.115 ;
    END
  END N4BEG[2]
  PIN N4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 32.750 222.315 33.030 223.115 ;
    END
  END N4BEG[3]
  PIN N4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 34.130 222.315 34.410 223.115 ;
    END
  END N4BEG[4]
  PIN N4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 35.510 222.315 35.790 223.115 ;
    END
  END N4BEG[5]
  PIN N4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 36.890 222.315 37.170 223.115 ;
    END
  END N4BEG[6]
  PIN N4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 38.270 222.315 38.550 223.115 ;
    END
  END N4BEG[7]
  PIN N4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 39.650 222.315 39.930 223.115 ;
    END
  END N4BEG[8]
  PIN N4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 41.030 222.315 41.310 223.115 ;
    END
  END N4BEG[9]
  PIN N4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 28.610 0.000 28.890 0.800 ;
    END
  END N4END[0]
  PIN N4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 42.410 0.000 42.690 0.800 ;
    END
  END N4END[10]
  PIN N4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 43.790 0.000 44.070 0.800 ;
    END
  END N4END[11]
  PIN N4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 0.800 ;
    END
  END N4END[12]
  PIN N4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 46.550 0.000 46.830 0.800 ;
    END
  END N4END[13]
  PIN N4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 47.930 0.000 48.210 0.800 ;
    END
  END N4END[14]
  PIN N4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 49.310 0.000 49.590 0.800 ;
    END
  END N4END[15]
  PIN N4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 29.990 0.000 30.270 0.800 ;
    END
  END N4END[1]
  PIN N4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 31.370 0.000 31.650 0.800 ;
    END
  END N4END[2]
  PIN N4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 32.750 0.000 33.030 0.800 ;
    END
  END N4END[3]
  PIN N4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 34.130 0.000 34.410 0.800 ;
    END
  END N4END[4]
  PIN N4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 0.800 ;
    END
  END N4END[5]
  PIN N4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 36.890 0.000 37.170 0.800 ;
    END
  END N4END[6]
  PIN N4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 38.270 0.000 38.550 0.800 ;
    END
  END N4END[7]
  PIN N4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 39.650 0.000 39.930 0.800 ;
    END
  END N4END[8]
  PIN N4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 41.030 0.000 41.310 0.800 ;
    END
  END N4END[9]
  PIN RAM2FAB_D0_I0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 129.200 35.400 130.000 36.000 ;
    END
  END RAM2FAB_D0_I0
  PIN RAM2FAB_D0_I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 129.200 38.120 130.000 38.720 ;
    END
  END RAM2FAB_D0_I1
  PIN RAM2FAB_D0_I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 129.200 40.840 130.000 41.440 ;
    END
  END RAM2FAB_D0_I2
  PIN RAM2FAB_D0_I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 129.200 43.560 130.000 44.160 ;
    END
  END RAM2FAB_D0_I3
  PIN RAM2FAB_D1_I0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 129.200 24.520 130.000 25.120 ;
    END
  END RAM2FAB_D1_I0
  PIN RAM2FAB_D1_I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 129.200 27.240 130.000 27.840 ;
    END
  END RAM2FAB_D1_I1
  PIN RAM2FAB_D1_I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 129.200 29.960 130.000 30.560 ;
    END
  END RAM2FAB_D1_I2
  PIN RAM2FAB_D1_I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 129.200 32.680 130.000 33.280 ;
    END
  END RAM2FAB_D1_I3
  PIN RAM2FAB_D2_I0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 129.200 13.640 130.000 14.240 ;
    END
  END RAM2FAB_D2_I0
  PIN RAM2FAB_D2_I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 129.200 16.360 130.000 16.960 ;
    END
  END RAM2FAB_D2_I1
  PIN RAM2FAB_D2_I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 129.200 19.080 130.000 19.680 ;
    END
  END RAM2FAB_D2_I2
  PIN RAM2FAB_D2_I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 129.200 21.800 130.000 22.400 ;
    END
  END RAM2FAB_D2_I3
  PIN RAM2FAB_D3_I0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 129.200 2.760 130.000 3.360 ;
    END
  END RAM2FAB_D3_I0
  PIN RAM2FAB_D3_I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 129.200 5.480 130.000 6.080 ;
    END
  END RAM2FAB_D3_I1
  PIN RAM2FAB_D3_I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 129.200 8.200 130.000 8.800 ;
    END
  END RAM2FAB_D3_I2
  PIN RAM2FAB_D3_I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 129.200 10.920 130.000 11.520 ;
    END
  END RAM2FAB_D3_I3
  PIN S1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 50.690 0.000 50.970 0.800 ;
    END
  END S1BEG[0]
  PIN S1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 52.070 0.000 52.350 0.800 ;
    END
  END S1BEG[1]
  PIN S1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 53.450 0.000 53.730 0.800 ;
    END
  END S1BEG[2]
  PIN S1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 0.800 ;
    END
  END S1BEG[3]
  PIN S1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 50.690 222.315 50.970 223.115 ;
    END
  END S1END[0]
  PIN S1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 52.070 222.315 52.350 223.115 ;
    END
  END S1END[1]
  PIN S1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 53.450 222.315 53.730 223.115 ;
    END
  END S1END[2]
  PIN S1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 54.830 222.315 55.110 223.115 ;
    END
  END S1END[3]
  PIN S2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 67.250 0.000 67.530 0.800 ;
    END
  END S2BEG[0]
  PIN S2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 68.630 0.000 68.910 0.800 ;
    END
  END S2BEG[1]
  PIN S2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 70.010 0.000 70.290 0.800 ;
    END
  END S2BEG[2]
  PIN S2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 71.390 0.000 71.670 0.800 ;
    END
  END S2BEG[3]
  PIN S2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 72.770 0.000 73.050 0.800 ;
    END
  END S2BEG[4]
  PIN S2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 0.800 ;
    END
  END S2BEG[5]
  PIN S2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 75.530 0.000 75.810 0.800 ;
    END
  END S2BEG[6]
  PIN S2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 76.910 0.000 77.190 0.800 ;
    END
  END S2BEG[7]
  PIN S2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 56.210 0.000 56.490 0.800 ;
    END
  END S2BEGb[0]
  PIN S2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 57.590 0.000 57.870 0.800 ;
    END
  END S2BEGb[1]
  PIN S2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 58.970 0.000 59.250 0.800 ;
    END
  END S2BEGb[2]
  PIN S2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 60.350 0.000 60.630 0.800 ;
    END
  END S2BEGb[3]
  PIN S2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 61.730 0.000 62.010 0.800 ;
    END
  END S2BEGb[4]
  PIN S2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 63.110 0.000 63.390 0.800 ;
    END
  END S2BEGb[5]
  PIN S2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 0.800 ;
    END
  END S2BEGb[6]
  PIN S2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 65.870 0.000 66.150 0.800 ;
    END
  END S2BEGb[7]
  PIN S2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 56.210 222.315 56.490 223.115 ;
    END
  END S2END[0]
  PIN S2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 57.590 222.315 57.870 223.115 ;
    END
  END S2END[1]
  PIN S2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 58.970 222.315 59.250 223.115 ;
    END
  END S2END[2]
  PIN S2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 60.350 222.315 60.630 223.115 ;
    END
  END S2END[3]
  PIN S2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 61.730 222.315 62.010 223.115 ;
    END
  END S2END[4]
  PIN S2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 63.110 222.315 63.390 223.115 ;
    END
  END S2END[5]
  PIN S2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 64.490 222.315 64.770 223.115 ;
    END
  END S2END[6]
  PIN S2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 65.870 222.315 66.150 223.115 ;
    END
  END S2END[7]
  PIN S2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 67.250 222.315 67.530 223.115 ;
    END
  END S2MID[0]
  PIN S2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 68.630 222.315 68.910 223.115 ;
    END
  END S2MID[1]
  PIN S2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 70.010 222.315 70.290 223.115 ;
    END
  END S2MID[2]
  PIN S2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 71.390 222.315 71.670 223.115 ;
    END
  END S2MID[3]
  PIN S2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 72.770 222.315 73.050 223.115 ;
    END
  END S2MID[4]
  PIN S2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 74.150 222.315 74.430 223.115 ;
    END
  END S2MID[5]
  PIN S2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 75.530 222.315 75.810 223.115 ;
    END
  END S2MID[6]
  PIN S2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 76.910 222.315 77.190 223.115 ;
    END
  END S2MID[7]
  PIN S4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 78.290 0.000 78.570 0.800 ;
    END
  END S4BEG[0]
  PIN S4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 92.090 0.000 92.370 0.800 ;
    END
  END S4BEG[10]
  PIN S4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 0.800 ;
    END
  END S4BEG[11]
  PIN S4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 94.850 0.000 95.130 0.800 ;
    END
  END S4BEG[12]
  PIN S4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 96.230 0.000 96.510 0.800 ;
    END
  END S4BEG[13]
  PIN S4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 97.610 0.000 97.890 0.800 ;
    END
  END S4BEG[14]
  PIN S4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 98.990 0.000 99.270 0.800 ;
    END
  END S4BEG[15]
  PIN S4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 79.670 0.000 79.950 0.800 ;
    END
  END S4BEG[1]
  PIN S4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 81.050 0.000 81.330 0.800 ;
    END
  END S4BEG[2]
  PIN S4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 82.430 0.000 82.710 0.800 ;
    END
  END S4BEG[3]
  PIN S4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 0.800 ;
    END
  END S4BEG[4]
  PIN S4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 85.190 0.000 85.470 0.800 ;
    END
  END S4BEG[5]
  PIN S4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 86.570 0.000 86.850 0.800 ;
    END
  END S4BEG[6]
  PIN S4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 87.950 0.000 88.230 0.800 ;
    END
  END S4BEG[7]
  PIN S4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 89.330 0.000 89.610 0.800 ;
    END
  END S4BEG[8]
  PIN S4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 90.710 0.000 90.990 0.800 ;
    END
  END S4BEG[9]
  PIN S4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 78.290 222.315 78.570 223.115 ;
    END
  END S4END[0]
  PIN S4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 92.090 222.315 92.370 223.115 ;
    END
  END S4END[10]
  PIN S4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 93.470 222.315 93.750 223.115 ;
    END
  END S4END[11]
  PIN S4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 94.850 222.315 95.130 223.115 ;
    END
  END S4END[12]
  PIN S4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 96.230 222.315 96.510 223.115 ;
    END
  END S4END[13]
  PIN S4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 97.610 222.315 97.890 223.115 ;
    END
  END S4END[14]
  PIN S4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 98.990 222.315 99.270 223.115 ;
    END
  END S4END[15]
  PIN S4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 79.670 222.315 79.950 223.115 ;
    END
  END S4END[1]
  PIN S4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 81.050 222.315 81.330 223.115 ;
    END
  END S4END[2]
  PIN S4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 82.430 222.315 82.710 223.115 ;
    END
  END S4END[3]
  PIN S4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 83.810 222.315 84.090 223.115 ;
    END
  END S4END[4]
  PIN S4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 85.190 222.315 85.470 223.115 ;
    END
  END S4END[5]
  PIN S4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 86.570 222.315 86.850 223.115 ;
    END
  END S4END[6]
  PIN S4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 87.950 222.315 88.230 223.115 ;
    END
  END S4END[7]
  PIN S4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 89.330 222.315 89.610 223.115 ;
    END
  END S4END[8]
  PIN S4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 90.710 222.315 90.990 223.115 ;
    END
  END S4END[9]
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 7.848000 ;
    PORT
      LAYER met2 ;
        RECT 100.370 0.000 100.650 0.800 ;
    END
  END UserCLK
  PIN UserCLKo
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 100.370 222.315 100.650 223.115 ;
    END
  END UserCLKo
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 34.390 5.200 35.990 217.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 64.060 5.200 65.660 217.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 93.730 5.200 95.330 217.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 123.400 5.200 125.000 217.840 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 19.555 5.200 21.155 217.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 49.225 5.200 50.825 217.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.895 5.200 80.495 217.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 108.565 5.200 110.165 217.840 ;
    END
  END VPWR
  PIN W1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 0.800 25.120 ;
    END
  END W1BEG[0]
  PIN W1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 0.800 26.480 ;
    END
  END W1BEG[1]
  PIN W1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 0.800 27.840 ;
    END
  END W1BEG[2]
  PIN W1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 0.800 29.200 ;
    END
  END W1BEG[3]
  PIN W2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 0.800 30.560 ;
    END
  END W2BEG[0]
  PIN W2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 0.800 31.920 ;
    END
  END W2BEG[1]
  PIN W2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 0.800 33.280 ;
    END
  END W2BEG[2]
  PIN W2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 0.800 34.640 ;
    END
  END W2BEG[3]
  PIN W2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 0.800 36.000 ;
    END
  END W2BEG[4]
  PIN W2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.760 0.800 37.360 ;
    END
  END W2BEG[5]
  PIN W2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 0.800 38.720 ;
    END
  END W2BEG[6]
  PIN W2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 0.800 40.080 ;
    END
  END W2BEG[7]
  PIN W2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 0.800 41.440 ;
    END
  END W2BEGb[0]
  PIN W2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 0.800 42.800 ;
    END
  END W2BEGb[1]
  PIN W2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 0.800 44.160 ;
    END
  END W2BEGb[2]
  PIN W2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 0.800 45.520 ;
    END
  END W2BEGb[3]
  PIN W2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 0.800 46.880 ;
    END
  END W2BEGb[4]
  PIN W2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 0.800 48.240 ;
    END
  END W2BEGb[5]
  PIN W2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 0.800 49.600 ;
    END
  END W2BEGb[6]
  PIN W2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 0.800 50.960 ;
    END
  END W2BEGb[7]
  PIN W6BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.480 0.800 74.080 ;
    END
  END W6BEG[0]
  PIN W6BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 0.800 87.680 ;
    END
  END W6BEG[10]
  PIN W6BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 0.800 89.040 ;
    END
  END W6BEG[11]
  PIN W6BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 0.800 75.440 ;
    END
  END W6BEG[1]
  PIN W6BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 0.800 76.800 ;
    END
  END W6BEG[2]
  PIN W6BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.560 0.800 78.160 ;
    END
  END W6BEG[3]
  PIN W6BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 0.800 79.520 ;
    END
  END W6BEG[4]
  PIN W6BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 0.800 80.880 ;
    END
  END W6BEG[5]
  PIN W6BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 0.800 82.240 ;
    END
  END W6BEG[6]
  PIN W6BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 0.800 83.600 ;
    END
  END W6BEG[7]
  PIN W6BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 0.800 84.960 ;
    END
  END W6BEG[8]
  PIN W6BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 0.800 86.320 ;
    END
  END W6BEG[9]
  PIN WW4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 0.800 52.320 ;
    END
  END WW4BEG[0]
  PIN WW4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 0.800 65.920 ;
    END
  END WW4BEG[10]
  PIN WW4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.680 0.800 67.280 ;
    END
  END WW4BEG[11]
  PIN WW4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 0.800 68.640 ;
    END
  END WW4BEG[12]
  PIN WW4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 0.800 70.000 ;
    END
  END WW4BEG[13]
  PIN WW4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 0.800 71.360 ;
    END
  END WW4BEG[14]
  PIN WW4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 0.800 72.720 ;
    END
  END WW4BEG[15]
  PIN WW4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 0.800 53.680 ;
    END
  END WW4BEG[1]
  PIN WW4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 0.800 55.040 ;
    END
  END WW4BEG[2]
  PIN WW4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 0.800 56.400 ;
    END
  END WW4BEG[3]
  PIN WW4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 0.800 57.760 ;
    END
  END WW4BEG[4]
  PIN WW4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 0.800 59.120 ;
    END
  END WW4BEG[5]
  PIN WW4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 0.800 60.480 ;
    END
  END WW4BEG[6]
  PIN WW4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 0.800 61.840 ;
    END
  END WW4BEG[7]
  PIN WW4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 0.800 63.200 ;
    END
  END WW4BEG[8]
  PIN WW4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 0.800 64.560 ;
    END
  END WW4BEG[9]
  OBS
      LAYER li1 ;
        RECT 5.520 5.355 124.200 217.685 ;
      LAYER met1 ;
        RECT 0.070 0.380 129.650 219.260 ;
      LAYER met2 ;
        RECT 0.100 222.035 0.730 222.315 ;
        RECT 1.570 222.035 2.110 222.315 ;
        RECT 2.950 222.035 3.490 222.315 ;
        RECT 4.330 222.035 4.870 222.315 ;
        RECT 5.710 222.035 6.250 222.315 ;
        RECT 7.090 222.035 7.630 222.315 ;
        RECT 8.470 222.035 9.010 222.315 ;
        RECT 9.850 222.035 10.390 222.315 ;
        RECT 11.230 222.035 11.770 222.315 ;
        RECT 12.610 222.035 13.150 222.315 ;
        RECT 13.990 222.035 14.530 222.315 ;
        RECT 15.370 222.035 15.910 222.315 ;
        RECT 16.750 222.035 17.290 222.315 ;
        RECT 18.130 222.035 18.670 222.315 ;
        RECT 19.510 222.035 20.050 222.315 ;
        RECT 20.890 222.035 21.430 222.315 ;
        RECT 22.270 222.035 22.810 222.315 ;
        RECT 23.650 222.035 24.190 222.315 ;
        RECT 25.030 222.035 25.570 222.315 ;
        RECT 26.410 222.035 26.950 222.315 ;
        RECT 27.790 222.035 28.330 222.315 ;
        RECT 29.170 222.035 29.710 222.315 ;
        RECT 30.550 222.035 31.090 222.315 ;
        RECT 31.930 222.035 32.470 222.315 ;
        RECT 33.310 222.035 33.850 222.315 ;
        RECT 34.690 222.035 35.230 222.315 ;
        RECT 36.070 222.035 36.610 222.315 ;
        RECT 37.450 222.035 37.990 222.315 ;
        RECT 38.830 222.035 39.370 222.315 ;
        RECT 40.210 222.035 40.750 222.315 ;
        RECT 41.590 222.035 42.130 222.315 ;
        RECT 42.970 222.035 43.510 222.315 ;
        RECT 44.350 222.035 44.890 222.315 ;
        RECT 45.730 222.035 46.270 222.315 ;
        RECT 47.110 222.035 47.650 222.315 ;
        RECT 48.490 222.035 49.030 222.315 ;
        RECT 49.870 222.035 50.410 222.315 ;
        RECT 51.250 222.035 51.790 222.315 ;
        RECT 52.630 222.035 53.170 222.315 ;
        RECT 54.010 222.035 54.550 222.315 ;
        RECT 55.390 222.035 55.930 222.315 ;
        RECT 56.770 222.035 57.310 222.315 ;
        RECT 58.150 222.035 58.690 222.315 ;
        RECT 59.530 222.035 60.070 222.315 ;
        RECT 60.910 222.035 61.450 222.315 ;
        RECT 62.290 222.035 62.830 222.315 ;
        RECT 63.670 222.035 64.210 222.315 ;
        RECT 65.050 222.035 65.590 222.315 ;
        RECT 66.430 222.035 66.970 222.315 ;
        RECT 67.810 222.035 68.350 222.315 ;
        RECT 69.190 222.035 69.730 222.315 ;
        RECT 70.570 222.035 71.110 222.315 ;
        RECT 71.950 222.035 72.490 222.315 ;
        RECT 73.330 222.035 73.870 222.315 ;
        RECT 74.710 222.035 75.250 222.315 ;
        RECT 76.090 222.035 76.630 222.315 ;
        RECT 77.470 222.035 78.010 222.315 ;
        RECT 78.850 222.035 79.390 222.315 ;
        RECT 80.230 222.035 80.770 222.315 ;
        RECT 81.610 222.035 82.150 222.315 ;
        RECT 82.990 222.035 83.530 222.315 ;
        RECT 84.370 222.035 84.910 222.315 ;
        RECT 85.750 222.035 86.290 222.315 ;
        RECT 87.130 222.035 87.670 222.315 ;
        RECT 88.510 222.035 89.050 222.315 ;
        RECT 89.890 222.035 90.430 222.315 ;
        RECT 91.270 222.035 91.810 222.315 ;
        RECT 92.650 222.035 93.190 222.315 ;
        RECT 94.030 222.035 94.570 222.315 ;
        RECT 95.410 222.035 95.950 222.315 ;
        RECT 96.790 222.035 97.330 222.315 ;
        RECT 98.170 222.035 98.710 222.315 ;
        RECT 99.550 222.035 100.090 222.315 ;
        RECT 100.930 222.035 101.470 222.315 ;
        RECT 102.310 222.035 102.850 222.315 ;
        RECT 103.690 222.035 104.230 222.315 ;
        RECT 105.070 222.035 105.610 222.315 ;
        RECT 106.450 222.035 106.990 222.315 ;
        RECT 107.830 222.035 108.370 222.315 ;
        RECT 109.210 222.035 109.750 222.315 ;
        RECT 110.590 222.035 111.130 222.315 ;
        RECT 111.970 222.035 112.510 222.315 ;
        RECT 113.350 222.035 113.890 222.315 ;
        RECT 114.730 222.035 115.270 222.315 ;
        RECT 116.110 222.035 116.650 222.315 ;
        RECT 117.490 222.035 118.030 222.315 ;
        RECT 118.870 222.035 119.410 222.315 ;
        RECT 120.250 222.035 120.790 222.315 ;
        RECT 121.630 222.035 122.170 222.315 ;
        RECT 123.010 222.035 123.550 222.315 ;
        RECT 124.390 222.035 124.930 222.315 ;
        RECT 125.770 222.035 126.310 222.315 ;
        RECT 127.150 222.035 127.690 222.315 ;
        RECT 128.530 222.035 129.630 222.315 ;
        RECT 0.100 1.080 129.630 222.035 ;
        RECT 0.100 0.270 0.730 1.080 ;
        RECT 1.570 0.270 2.110 1.080 ;
        RECT 2.950 0.270 3.490 1.080 ;
        RECT 4.330 0.270 4.870 1.080 ;
        RECT 5.710 0.270 6.250 1.080 ;
        RECT 7.090 0.270 7.630 1.080 ;
        RECT 8.470 0.270 9.010 1.080 ;
        RECT 9.850 0.270 10.390 1.080 ;
        RECT 11.230 0.270 11.770 1.080 ;
        RECT 12.610 0.270 13.150 1.080 ;
        RECT 13.990 0.270 14.530 1.080 ;
        RECT 15.370 0.270 15.910 1.080 ;
        RECT 16.750 0.270 17.290 1.080 ;
        RECT 18.130 0.270 18.670 1.080 ;
        RECT 19.510 0.270 20.050 1.080 ;
        RECT 20.890 0.270 21.430 1.080 ;
        RECT 22.270 0.270 22.810 1.080 ;
        RECT 23.650 0.270 24.190 1.080 ;
        RECT 25.030 0.270 25.570 1.080 ;
        RECT 26.410 0.270 26.950 1.080 ;
        RECT 27.790 0.270 28.330 1.080 ;
        RECT 29.170 0.270 29.710 1.080 ;
        RECT 30.550 0.270 31.090 1.080 ;
        RECT 31.930 0.270 32.470 1.080 ;
        RECT 33.310 0.270 33.850 1.080 ;
        RECT 34.690 0.270 35.230 1.080 ;
        RECT 36.070 0.270 36.610 1.080 ;
        RECT 37.450 0.270 37.990 1.080 ;
        RECT 38.830 0.270 39.370 1.080 ;
        RECT 40.210 0.270 40.750 1.080 ;
        RECT 41.590 0.270 42.130 1.080 ;
        RECT 42.970 0.270 43.510 1.080 ;
        RECT 44.350 0.270 44.890 1.080 ;
        RECT 45.730 0.270 46.270 1.080 ;
        RECT 47.110 0.270 47.650 1.080 ;
        RECT 48.490 0.270 49.030 1.080 ;
        RECT 49.870 0.270 50.410 1.080 ;
        RECT 51.250 0.270 51.790 1.080 ;
        RECT 52.630 0.270 53.170 1.080 ;
        RECT 54.010 0.270 54.550 1.080 ;
        RECT 55.390 0.270 55.930 1.080 ;
        RECT 56.770 0.270 57.310 1.080 ;
        RECT 58.150 0.270 58.690 1.080 ;
        RECT 59.530 0.270 60.070 1.080 ;
        RECT 60.910 0.270 61.450 1.080 ;
        RECT 62.290 0.270 62.830 1.080 ;
        RECT 63.670 0.270 64.210 1.080 ;
        RECT 65.050 0.270 65.590 1.080 ;
        RECT 66.430 0.270 66.970 1.080 ;
        RECT 67.810 0.270 68.350 1.080 ;
        RECT 69.190 0.270 69.730 1.080 ;
        RECT 70.570 0.270 71.110 1.080 ;
        RECT 71.950 0.270 72.490 1.080 ;
        RECT 73.330 0.270 73.870 1.080 ;
        RECT 74.710 0.270 75.250 1.080 ;
        RECT 76.090 0.270 76.630 1.080 ;
        RECT 77.470 0.270 78.010 1.080 ;
        RECT 78.850 0.270 79.390 1.080 ;
        RECT 80.230 0.270 80.770 1.080 ;
        RECT 81.610 0.270 82.150 1.080 ;
        RECT 82.990 0.270 83.530 1.080 ;
        RECT 84.370 0.270 84.910 1.080 ;
        RECT 85.750 0.270 86.290 1.080 ;
        RECT 87.130 0.270 87.670 1.080 ;
        RECT 88.510 0.270 89.050 1.080 ;
        RECT 89.890 0.270 90.430 1.080 ;
        RECT 91.270 0.270 91.810 1.080 ;
        RECT 92.650 0.270 93.190 1.080 ;
        RECT 94.030 0.270 94.570 1.080 ;
        RECT 95.410 0.270 95.950 1.080 ;
        RECT 96.790 0.270 97.330 1.080 ;
        RECT 98.170 0.270 98.710 1.080 ;
        RECT 99.550 0.270 100.090 1.080 ;
        RECT 100.930 0.270 101.470 1.080 ;
        RECT 102.310 0.270 102.850 1.080 ;
        RECT 103.690 0.270 104.230 1.080 ;
        RECT 105.070 0.270 105.610 1.080 ;
        RECT 106.450 0.270 106.990 1.080 ;
        RECT 107.830 0.270 108.370 1.080 ;
        RECT 109.210 0.270 109.750 1.080 ;
        RECT 110.590 0.270 111.130 1.080 ;
        RECT 111.970 0.270 112.510 1.080 ;
        RECT 113.350 0.270 113.890 1.080 ;
        RECT 114.730 0.270 115.270 1.080 ;
        RECT 116.110 0.270 116.650 1.080 ;
        RECT 117.490 0.270 118.030 1.080 ;
        RECT 118.870 0.270 119.410 1.080 ;
        RECT 120.250 0.270 120.790 1.080 ;
        RECT 121.630 0.270 122.170 1.080 ;
        RECT 123.010 0.270 123.550 1.080 ;
        RECT 124.390 0.270 124.930 1.080 ;
        RECT 125.770 0.270 126.310 1.080 ;
        RECT 127.150 0.270 127.690 1.080 ;
        RECT 128.530 0.270 129.630 1.080 ;
      LAYER met3 ;
        RECT 0.800 217.240 128.800 218.090 ;
        RECT 0.800 215.920 129.655 217.240 ;
        RECT 0.800 214.520 128.800 215.920 ;
        RECT 0.800 213.200 129.655 214.520 ;
        RECT 0.800 211.800 128.800 213.200 ;
        RECT 0.800 210.480 129.655 211.800 ;
        RECT 0.800 209.080 128.800 210.480 ;
        RECT 0.800 207.760 129.655 209.080 ;
        RECT 0.800 206.360 128.800 207.760 ;
        RECT 0.800 205.040 129.655 206.360 ;
        RECT 0.800 203.640 128.800 205.040 ;
        RECT 0.800 202.320 129.655 203.640 ;
        RECT 0.800 200.920 128.800 202.320 ;
        RECT 0.800 199.600 129.655 200.920 ;
        RECT 0.800 198.240 128.800 199.600 ;
        RECT 1.200 198.200 128.800 198.240 ;
        RECT 1.200 196.880 129.655 198.200 ;
        RECT 1.200 195.480 128.800 196.880 ;
        RECT 1.200 194.160 129.655 195.480 ;
        RECT 1.200 192.760 128.800 194.160 ;
        RECT 1.200 191.440 129.655 192.760 ;
        RECT 1.200 190.040 128.800 191.440 ;
        RECT 1.200 188.720 129.655 190.040 ;
        RECT 1.200 187.320 128.800 188.720 ;
        RECT 1.200 186.000 129.655 187.320 ;
        RECT 1.200 184.600 128.800 186.000 ;
        RECT 1.200 183.280 129.655 184.600 ;
        RECT 1.200 181.880 128.800 183.280 ;
        RECT 1.200 180.560 129.655 181.880 ;
        RECT 1.200 179.160 128.800 180.560 ;
        RECT 1.200 177.840 129.655 179.160 ;
        RECT 1.200 176.440 128.800 177.840 ;
        RECT 1.200 175.120 129.655 176.440 ;
        RECT 1.200 173.720 128.800 175.120 ;
        RECT 1.200 172.400 129.655 173.720 ;
        RECT 1.200 171.000 128.800 172.400 ;
        RECT 1.200 169.680 129.655 171.000 ;
        RECT 1.200 168.280 128.800 169.680 ;
        RECT 1.200 166.960 129.655 168.280 ;
        RECT 1.200 165.560 128.800 166.960 ;
        RECT 1.200 164.240 129.655 165.560 ;
        RECT 1.200 162.840 128.800 164.240 ;
        RECT 1.200 161.520 129.655 162.840 ;
        RECT 1.200 160.120 128.800 161.520 ;
        RECT 1.200 158.800 129.655 160.120 ;
        RECT 1.200 157.400 128.800 158.800 ;
        RECT 1.200 156.080 129.655 157.400 ;
        RECT 1.200 154.680 128.800 156.080 ;
        RECT 1.200 153.360 129.655 154.680 ;
        RECT 1.200 151.960 128.800 153.360 ;
        RECT 1.200 150.640 129.655 151.960 ;
        RECT 1.200 149.240 128.800 150.640 ;
        RECT 1.200 147.920 129.655 149.240 ;
        RECT 1.200 146.520 128.800 147.920 ;
        RECT 1.200 145.200 129.655 146.520 ;
        RECT 1.200 143.800 128.800 145.200 ;
        RECT 1.200 142.480 129.655 143.800 ;
        RECT 1.200 141.080 128.800 142.480 ;
        RECT 1.200 139.760 129.655 141.080 ;
        RECT 1.200 138.360 128.800 139.760 ;
        RECT 1.200 137.040 129.655 138.360 ;
        RECT 1.200 135.640 128.800 137.040 ;
        RECT 1.200 134.320 129.655 135.640 ;
        RECT 1.200 132.920 128.800 134.320 ;
        RECT 1.200 131.600 129.655 132.920 ;
        RECT 1.200 130.200 128.800 131.600 ;
        RECT 1.200 128.880 129.655 130.200 ;
        RECT 1.200 127.480 128.800 128.880 ;
        RECT 1.200 126.160 129.655 127.480 ;
        RECT 1.200 124.760 128.800 126.160 ;
        RECT 1.200 123.440 129.655 124.760 ;
        RECT 1.200 122.040 128.800 123.440 ;
        RECT 1.200 120.720 129.655 122.040 ;
        RECT 1.200 119.320 128.800 120.720 ;
        RECT 1.200 118.000 129.655 119.320 ;
        RECT 1.200 116.600 128.800 118.000 ;
        RECT 1.200 115.280 129.655 116.600 ;
        RECT 1.200 113.880 128.800 115.280 ;
        RECT 1.200 112.560 129.655 113.880 ;
        RECT 1.200 111.160 128.800 112.560 ;
        RECT 1.200 109.840 129.655 111.160 ;
        RECT 1.200 108.440 128.800 109.840 ;
        RECT 1.200 107.120 129.655 108.440 ;
        RECT 1.200 105.720 128.800 107.120 ;
        RECT 1.200 104.400 129.655 105.720 ;
        RECT 1.200 103.000 128.800 104.400 ;
        RECT 1.200 101.680 129.655 103.000 ;
        RECT 1.200 100.280 128.800 101.680 ;
        RECT 1.200 98.960 129.655 100.280 ;
        RECT 1.200 97.560 128.800 98.960 ;
        RECT 1.200 96.240 129.655 97.560 ;
        RECT 1.200 94.840 128.800 96.240 ;
        RECT 1.200 93.520 129.655 94.840 ;
        RECT 1.200 92.120 128.800 93.520 ;
        RECT 1.200 90.800 129.655 92.120 ;
        RECT 1.200 89.400 128.800 90.800 ;
        RECT 1.200 88.080 129.655 89.400 ;
        RECT 1.200 86.680 128.800 88.080 ;
        RECT 1.200 85.360 129.655 86.680 ;
        RECT 1.200 83.960 128.800 85.360 ;
        RECT 1.200 82.640 129.655 83.960 ;
        RECT 1.200 81.240 128.800 82.640 ;
        RECT 1.200 79.920 129.655 81.240 ;
        RECT 1.200 78.520 128.800 79.920 ;
        RECT 1.200 77.200 129.655 78.520 ;
        RECT 1.200 75.800 128.800 77.200 ;
        RECT 1.200 74.480 129.655 75.800 ;
        RECT 1.200 73.080 128.800 74.480 ;
        RECT 1.200 71.760 129.655 73.080 ;
        RECT 1.200 70.360 128.800 71.760 ;
        RECT 1.200 69.040 129.655 70.360 ;
        RECT 1.200 67.640 128.800 69.040 ;
        RECT 1.200 66.320 129.655 67.640 ;
        RECT 1.200 64.920 128.800 66.320 ;
        RECT 1.200 63.600 129.655 64.920 ;
        RECT 1.200 62.200 128.800 63.600 ;
        RECT 1.200 60.880 129.655 62.200 ;
        RECT 1.200 59.480 128.800 60.880 ;
        RECT 1.200 58.160 129.655 59.480 ;
        RECT 1.200 56.760 128.800 58.160 ;
        RECT 1.200 55.440 129.655 56.760 ;
        RECT 1.200 54.040 128.800 55.440 ;
        RECT 1.200 52.720 129.655 54.040 ;
        RECT 1.200 51.320 128.800 52.720 ;
        RECT 1.200 50.000 129.655 51.320 ;
        RECT 1.200 48.600 128.800 50.000 ;
        RECT 1.200 47.280 129.655 48.600 ;
        RECT 1.200 45.880 128.800 47.280 ;
        RECT 1.200 44.560 129.655 45.880 ;
        RECT 1.200 43.160 128.800 44.560 ;
        RECT 1.200 41.840 129.655 43.160 ;
        RECT 1.200 40.440 128.800 41.840 ;
        RECT 1.200 39.120 129.655 40.440 ;
        RECT 1.200 37.720 128.800 39.120 ;
        RECT 1.200 36.400 129.655 37.720 ;
        RECT 1.200 35.000 128.800 36.400 ;
        RECT 1.200 33.680 129.655 35.000 ;
        RECT 1.200 32.280 128.800 33.680 ;
        RECT 1.200 30.960 129.655 32.280 ;
        RECT 1.200 29.560 128.800 30.960 ;
        RECT 1.200 28.240 129.655 29.560 ;
        RECT 1.200 26.840 128.800 28.240 ;
        RECT 1.200 25.520 129.655 26.840 ;
        RECT 1.200 24.120 128.800 25.520 ;
        RECT 0.800 22.800 129.655 24.120 ;
        RECT 0.800 21.400 128.800 22.800 ;
        RECT 0.800 20.080 129.655 21.400 ;
        RECT 0.800 18.680 128.800 20.080 ;
        RECT 0.800 17.360 129.655 18.680 ;
        RECT 0.800 15.960 128.800 17.360 ;
        RECT 0.800 14.640 129.655 15.960 ;
        RECT 0.800 13.240 128.800 14.640 ;
        RECT 0.800 11.920 129.655 13.240 ;
        RECT 0.800 10.520 128.800 11.920 ;
        RECT 0.800 9.200 129.655 10.520 ;
        RECT 0.800 7.800 128.800 9.200 ;
        RECT 0.800 6.480 129.655 7.800 ;
        RECT 0.800 5.080 128.800 6.480 ;
        RECT 0.800 3.760 129.655 5.080 ;
        RECT 0.800 2.895 128.800 3.760 ;
      LAYER met4 ;
        RECT 3.055 5.615 19.155 214.705 ;
        RECT 21.555 5.615 33.990 214.705 ;
        RECT 36.390 5.615 48.825 214.705 ;
        RECT 51.225 5.615 63.660 214.705 ;
        RECT 66.060 5.615 78.495 214.705 ;
        RECT 80.895 5.615 93.330 214.705 ;
        RECT 95.730 5.615 108.165 214.705 ;
        RECT 110.565 5.615 114.705 214.705 ;
  END
END RAM_IO
END LIBRARY

